// RTL (Verilog) generated @ Sun Feb 20 16:09:27 2022 by V3 
//               compiled @ Feb 20 2022 16:07:45
// Internal nets are renamed with prefix "v3_1645344567_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1645344567_0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] v3_1645344567_8;
   reg [2:0] v3_1645344567_9;
   reg [2:0] v3_1645344567_10;
   reg [2:0] v3_1645344567_11;
   reg [1:0] v3_1645344567_12;
   reg [1:0] v3_1645344567_13;
   reg v3_1645344567_14;
   reg [7:0] v3_1645344567_15;
   reg v3_1645344567_16;
   reg [1:0] v3_1645344567_17;
   reg [7:0] v3_1645344567_18;
   reg [2:0] v3_1645344567_19;
   reg [2:0] v3_1645344567_20;
   reg [2:0] v3_1645344567_21;
   reg [2:0] v3_1645344567_22;
   wire [2:0] v3_1645344567_23;
   wire [2:0] v3_1645344567_24;
   wire [2:0] v3_1645344567_25;
   wire [2:0] v3_1645344567_26;
   wire [2:0] v3_1645344567_27;
   wire [2:0] v3_1645344567_28;
   wire [2:0] v3_1645344567_29;
   wire [2:0] v3_1645344567_30;
   wire [2:0] v3_1645344567_31;
   wire [2:0] v3_1645344567_32;
   wire [2:0] v3_1645344567_33;
   wire [2:0] v3_1645344567_34;
   wire [2:0] v3_1645344567_35;
   wire v3_1645344567_36;
   wire v3_1645344567_37;
   wire [7:0] v3_1645344567_38;
   wire v3_1645344567_39;
   wire [1:0] v3_1645344567_40;
   wire v3_1645344567_41;
   wire [1:0] v3_1645344567_42;
   wire [2:0] v3_1645344567_43;
   wire [2:0] v3_1645344567_44;
   wire [2:0] v3_1645344567_45;
   wire [2:0] v3_1645344567_46;
   wire [2:0] v3_1645344567_47;
   wire v3_1645344567_48;
   wire v3_1645344567_49;
   wire [7:0] v3_1645344567_50;
   wire v3_1645344567_51;
   wire [1:0] v3_1645344567_52;
   wire v3_1645344567_53;
   wire [2:0] v3_1645344567_54;
   wire v3_1645344567_55;
   wire [2:0] v3_1645344567_56;
   wire [2:0] v3_1645344567_57;
   wire v3_1645344567_58;
   wire v3_1645344567_59;
   wire v3_1645344567_60;
   wire [2:0] v3_1645344567_61;
   wire v3_1645344567_62;
   wire [2:0] v3_1645344567_63;
   wire [2:0] v3_1645344567_64;
   wire [2:0] v3_1645344567_65;
   wire [2:0] v3_1645344567_66;
   wire [2:0] v3_1645344567_67;
   wire [2:0] v3_1645344567_68;
   wire [2:0] v3_1645344567_69;
   wire [2:0] v3_1645344567_70;
   wire [2:0] v3_1645344567_71;
   wire [2:0] v3_1645344567_72;
   wire [2:0] v3_1645344567_73;
   wire [2:0] v3_1645344567_74;
   wire [2:0] v3_1645344567_75;
   wire [2:0] v3_1645344567_76;
   wire [2:0] v3_1645344567_77;
   wire [2:0] v3_1645344567_78;
   wire [2:0] v3_1645344567_79;
   wire v3_1645344567_80;
   wire v3_1645344567_81;
   wire [7:0] v3_1645344567_82;
   wire [2:0] v3_1645344567_83;
   wire [2:0] v3_1645344567_84;
   wire [2:0] v3_1645344567_85;
   wire [2:0] v3_1645344567_86;
   wire [2:0] v3_1645344567_87;
   wire [2:0] v3_1645344567_88;
   wire [2:0] v3_1645344567_89;
   wire [2:0] v3_1645344567_90;
   wire [2:0] v3_1645344567_91;
   wire [2:0] v3_1645344567_92;
   wire [2:0] v3_1645344567_93;
   wire [2:0] v3_1645344567_94;
   wire [2:0] v3_1645344567_95;
   wire [2:0] v3_1645344567_96;
   wire [2:0] v3_1645344567_97;
   wire [2:0] v3_1645344567_98;
   wire [2:0] v3_1645344567_99;
   wire [2:0] v3_1645344567_100;
   wire [2:0] v3_1645344567_101;
   wire [2:0] v3_1645344567_102;
   wire [2:0] v3_1645344567_103;
   wire v3_1645344567_104;
   wire v3_1645344567_105;
   wire [7:0] v3_1645344567_106;
   wire [2:0] v3_1645344567_107;
   wire [2:0] v3_1645344567_108;
   wire [2:0] v3_1645344567_109;
   wire [2:0] v3_1645344567_110;
   wire [2:0] v3_1645344567_111;
   wire [2:0] v3_1645344567_112;
   wire [2:0] v3_1645344567_113;
   wire [2:0] v3_1645344567_114;
   wire [2:0] v3_1645344567_115;
   wire [2:0] v3_1645344567_116;
   wire [2:0] v3_1645344567_117;
   wire [2:0] v3_1645344567_118;
   wire [2:0] v3_1645344567_119;
   wire [2:0] v3_1645344567_120;
   wire [2:0] v3_1645344567_121;
   wire [2:0] v3_1645344567_122;
   wire [2:0] v3_1645344567_123;
   wire [2:0] v3_1645344567_124;
   wire [2:0] v3_1645344567_125;
   wire [2:0] v3_1645344567_126;
   wire [2:0] v3_1645344567_127;
   wire [2:0] v3_1645344567_128;
   wire [2:0] v3_1645344567_129;
   wire [2:0] v3_1645344567_130;
   wire [1:0] v3_1645344567_131;
   wire [1:0] v3_1645344567_132;
   wire [1:0] v3_1645344567_133;
   wire [1:0] v3_1645344567_134;
   wire [1:0] v3_1645344567_135;
   wire [1:0] v3_1645344567_136;
   wire [1:0] v3_1645344567_137;
   wire [1:0] v3_1645344567_138;
   wire [1:0] v3_1645344567_139;
   wire [1:0] v3_1645344567_140;
   wire [1:0] v3_1645344567_141;
   wire [1:0] v3_1645344567_142;
   wire [1:0] v3_1645344567_143;
   wire [1:0] v3_1645344567_144;
   wire v3_1645344567_145;
   wire v3_1645344567_146;
   wire [1:0] v3_1645344567_147;
   wire [1:0] v3_1645344567_148;
   wire [1:0] v3_1645344567_149;
   wire [1:0] v3_1645344567_150;
   wire [1:0] v3_1645344567_151;
   wire [1:0] v3_1645344567_152;
   wire [1:0] v3_1645344567_153;
   wire [1:0] v3_1645344567_154;
   wire [1:0] v3_1645344567_155;
   wire [1:0] v3_1645344567_156;
   wire [1:0] v3_1645344567_157;
   wire [1:0] v3_1645344567_158;
   wire [1:0] v3_1645344567_159;
   wire [1:0] v3_1645344567_160;
   wire [1:0] v3_1645344567_161;
   wire [1:0] v3_1645344567_162;
   wire [1:0] v3_1645344567_163;
   wire [1:0] v3_1645344567_164;
   wire [1:0] v3_1645344567_165;
   wire [1:0] v3_1645344567_166;
   wire [1:0] v3_1645344567_167;
   wire [1:0] v3_1645344567_168;
   wire [1:0] v3_1645344567_169;
   wire v3_1645344567_170;
   wire v3_1645344567_171;
   wire v3_1645344567_172;
   wire v3_1645344567_173;
   wire v3_1645344567_174;
   wire [7:0] v3_1645344567_175;
   wire [7:0] v3_1645344567_176;
   wire [7:0] v3_1645344567_177;
   wire [7:0] v3_1645344567_178;
   wire [7:0] v3_1645344567_179;
   wire [7:0] v3_1645344567_180;
   wire [7:0] v3_1645344567_181;
   wire [7:0] v3_1645344567_182;
   wire [7:0] v3_1645344567_183;
   wire [7:0] v3_1645344567_184;
   wire [5:0] v3_1645344567_185;
   wire [7:0] v3_1645344567_186;
   wire [7:0] v3_1645344567_187;
   wire [7:0] v3_1645344567_188;
   wire [7:0] v3_1645344567_189;
   wire [7:0] v3_1645344567_190;
   wire [7:0] v3_1645344567_191;
   wire [7:0] v3_1645344567_192;
   wire [7:0] v3_1645344567_193;
   wire [7:0] v3_1645344567_194;
   wire [7:0] v3_1645344567_195;
   wire [7:0] v3_1645344567_196;
   wire [7:0] v3_1645344567_197;
   wire [7:0] v3_1645344567_198;
   wire [7:0] v3_1645344567_199;
   wire [7:0] v3_1645344567_200;
   wire [7:0] v3_1645344567_201;
   wire [7:0] v3_1645344567_202;
   wire [7:0] v3_1645344567_203;
   wire [7:0] v3_1645344567_204;
   wire [7:0] v3_1645344567_205;
   wire v3_1645344567_206;
   wire v3_1645344567_207;
   wire v3_1645344567_208;
   wire v3_1645344567_209;
   wire v3_1645344567_210;
   wire v3_1645344567_211;
   wire v3_1645344567_212;
   wire v3_1645344567_213;
   wire v3_1645344567_214;
   wire v3_1645344567_215;
   wire v3_1645344567_216;
   wire v3_1645344567_217;
   wire v3_1645344567_218;
   wire v3_1645344567_219;
   wire [1:0] v3_1645344567_220;
   wire [1:0] v3_1645344567_221;
   wire [1:0] v3_1645344567_222;
   wire [1:0] v3_1645344567_223;
   wire [1:0] v3_1645344567_224;
   wire [1:0] v3_1645344567_225;
   wire [1:0] v3_1645344567_226;
   wire [1:0] v3_1645344567_227;
   wire [1:0] v3_1645344567_228;
   wire [1:0] v3_1645344567_229;
   wire [1:0] v3_1645344567_230;
   wire [1:0] v3_1645344567_231;
   wire [1:0] v3_1645344567_232;
   wire [1:0] v3_1645344567_233;
   wire [1:0] v3_1645344567_234;
   wire [1:0] v3_1645344567_235;
   wire [1:0] v3_1645344567_236;
   wire [1:0] v3_1645344567_237;
   wire [1:0] v3_1645344567_238;
   wire [1:0] v3_1645344567_239;
   wire [1:0] v3_1645344567_240;
   wire [1:0] v3_1645344567_241;
   wire [1:0] v3_1645344567_242;
   wire [1:0] v3_1645344567_243;
   wire [1:0] v3_1645344567_244;
   wire [1:0] v3_1645344567_245;
   wire [1:0] v3_1645344567_246;
   wire [1:0] v3_1645344567_247;
   wire [1:0] v3_1645344567_248;
   wire [7:0] v3_1645344567_249;
   wire [7:0] v3_1645344567_250;
   wire [7:0] v3_1645344567_251;
   wire [7:0] v3_1645344567_252;
   wire [7:0] v3_1645344567_253;
   wire [7:0] v3_1645344567_254;
   wire [7:0] v3_1645344567_255;
   wire [7:0] v3_1645344567_256;
   wire [7:0] v3_1645344567_257;
   wire [7:0] v3_1645344567_258;
   wire [7:0] v3_1645344567_259;
   wire [7:0] v3_1645344567_260;
   wire [7:0] v3_1645344567_261;
   wire [7:0] v3_1645344567_262;
   wire [7:0] v3_1645344567_263;
   wire [7:0] v3_1645344567_264;
   wire [7:0] v3_1645344567_265;
   wire [7:0] v3_1645344567_266;
   wire [7:0] v3_1645344567_267;
   wire [7:0] v3_1645344567_268;
   wire [7:0] v3_1645344567_269;
   wire [7:0] v3_1645344567_270;
   wire [7:0] v3_1645344567_271;
   wire [7:0] v3_1645344567_272;
   wire [7:0] v3_1645344567_273;
   wire [7:0] v3_1645344567_274;
   wire [7:0] v3_1645344567_275;
   wire [7:0] v3_1645344567_276;
   wire [7:0] v3_1645344567_277;
   wire [7:0] v3_1645344567_278;
   wire [7:0] v3_1645344567_279;
   wire [7:0] v3_1645344567_280;
   wire [7:0] v3_1645344567_281;
   wire [7:0] v3_1645344567_282;
   wire [7:0] v3_1645344567_283;
   wire v3_1645344567_284;
   wire [7:0] v3_1645344567_285;
   wire v3_1645344567_286;
   wire [7:0] v3_1645344567_287;
   wire v3_1645344567_288;
   wire [7:0] v3_1645344567_289;
   wire [7:0] v3_1645344567_290;
   wire [2:0] v3_1645344567_291;
   wire [2:0] v3_1645344567_292;
   wire [2:0] v3_1645344567_293;
   wire [2:0] v3_1645344567_294;
   wire [2:0] v3_1645344567_295;
   wire [2:0] v3_1645344567_296;
   wire [2:0] v3_1645344567_297;
   wire [2:0] v3_1645344567_298;
   wire [2:0] v3_1645344567_299;
   wire [2:0] v3_1645344567_300;
   wire [2:0] v3_1645344567_301;
   wire [2:0] v3_1645344567_302;
   wire [2:0] v3_1645344567_303;
   wire [2:0] v3_1645344567_304;
   wire [2:0] v3_1645344567_305;
   wire [2:0] v3_1645344567_306;
   wire [2:0] v3_1645344567_307;
   wire [2:0] v3_1645344567_308;
   wire [2:0] v3_1645344567_309;
   wire [2:0] v3_1645344567_310;
   wire [2:0] v3_1645344567_311;
   wire [2:0] v3_1645344567_312;
   wire [2:0] v3_1645344567_313;
   wire [2:0] v3_1645344567_314;
   wire v3_1645344567_315;
   wire [3:0] v3_1645344567_316;
   wire [3:0] v3_1645344567_317;
   wire [3:0] v3_1645344567_318;
   wire [3:0] v3_1645344567_319;
   wire [3:0] v3_1645344567_320;
   wire [3:0] v3_1645344567_321;
   wire [3:0] v3_1645344567_322;
   wire [2:0] v3_1645344567_323;
   wire [2:0] v3_1645344567_324;
   wire [2:0] v3_1645344567_325;
   wire [2:0] v3_1645344567_326;
   wire [2:0] v3_1645344567_327;
   wire [2:0] v3_1645344567_328;
   wire [2:0] v3_1645344567_329;
   wire [2:0] v3_1645344567_330;
   wire [2:0] v3_1645344567_331;
   wire [2:0] v3_1645344567_332;
   wire [2:0] v3_1645344567_333;
   wire [2:0] v3_1645344567_334;
   wire [2:0] v3_1645344567_335;
   wire [2:0] v3_1645344567_336;
   wire [2:0] v3_1645344567_337;
   wire [2:0] v3_1645344567_338;
   wire [2:0] v3_1645344567_339;
   wire [2:0] v3_1645344567_340;
   wire [2:0] v3_1645344567_341;
   wire [2:0] v3_1645344567_342;
   wire [2:0] v3_1645344567_343;
   wire [2:0] v3_1645344567_344;
   wire [2:0] v3_1645344567_345;
   wire [2:0] v3_1645344567_346;
   wire [2:0] v3_1645344567_347;
   wire [2:0] v3_1645344567_348;
   wire v3_1645344567_349;
   wire [3:0] v3_1645344567_350;
   wire [3:0] v3_1645344567_351;
   wire [3:0] v3_1645344567_352;
   wire [3:0] v3_1645344567_353;
   wire [3:0] v3_1645344567_354;
   wire [3:0] v3_1645344567_355;
   wire [2:0] v3_1645344567_356;
   wire [2:0] v3_1645344567_357;
   wire [2:0] v3_1645344567_358;
   wire [2:0] v3_1645344567_359;
   wire [2:0] v3_1645344567_360;
   wire [2:0] v3_1645344567_361;
   wire [2:0] v3_1645344567_362;
   wire [2:0] v3_1645344567_363;
   wire [2:0] v3_1645344567_364;
   wire [2:0] v3_1645344567_365;
   wire [2:0] v3_1645344567_366;
   wire [2:0] v3_1645344567_367;
   wire [2:0] v3_1645344567_368;
   wire [2:0] v3_1645344567_369;
   wire [2:0] v3_1645344567_370;
   wire [2:0] v3_1645344567_371;
   wire [2:0] v3_1645344567_372;
   wire [2:0] v3_1645344567_373;
   wire [2:0] v3_1645344567_374;
   wire [2:0] v3_1645344567_375;
   wire [2:0] v3_1645344567_376;
   wire [2:0] v3_1645344567_377;
   wire [2:0] v3_1645344567_378;
   wire v3_1645344567_379;
   wire [3:0] v3_1645344567_380;
   wire [3:0] v3_1645344567_381;
   wire [3:0] v3_1645344567_382;
   wire [3:0] v3_1645344567_383;
   wire [3:0] v3_1645344567_384;
   wire [3:0] v3_1645344567_385;
   wire [2:0] v3_1645344567_386;
   wire [2:0] v3_1645344567_387;
   wire [2:0] v3_1645344567_388;
   wire [2:0] v3_1645344567_389;
   wire [2:0] v3_1645344567_390;
   wire [2:0] v3_1645344567_391;
   wire [2:0] v3_1645344567_392;
   wire [2:0] v3_1645344567_393;
   wire [2:0] v3_1645344567_394;
   wire [2:0] v3_1645344567_395;
   wire [2:0] v3_1645344567_396;
   wire [2:0] v3_1645344567_397;
   wire [2:0] v3_1645344567_398;
   wire [2:0] v3_1645344567_399;
   wire [2:0] v3_1645344567_400;
   wire [2:0] v3_1645344567_401;
   wire [2:0] v3_1645344567_402;
   wire [2:0] v3_1645344567_403;
   wire [2:0] v3_1645344567_404;
   wire [2:0] v3_1645344567_405;
   wire [2:0] v3_1645344567_406;
   wire [2:0] v3_1645344567_407;
   wire [2:0] v3_1645344567_408;
   wire [2:0] v3_1645344567_409;
   wire [2:0] v3_1645344567_410;
   wire v3_1645344567_411;
   wire [3:0] v3_1645344567_412;
   wire [3:0] v3_1645344567_413;
   wire [3:0] v3_1645344567_414;
   wire [3:0] v3_1645344567_415;
   wire [3:0] v3_1645344567_416;
   wire [3:0] v3_1645344567_417;
   wire [2:0] v3_1645344567_418;
   wire [2:0] v3_1645344567_419;
   wire v3_1645344567_420;
   wire v3_1645344567_421;
   wire v3_1645344567_422;
   wire v3_1645344567_423;
   wire v3_1645344567_424;
   wire v3_1645344567_425;
   wire v3_1645344567_426;
   wire v3_1645344567_427;
   wire [7:0] v3_1645344567_428;
   wire [7:0] v3_1645344567_429;
   wire [7:0] v3_1645344567_430;
   wire [7:0] v3_1645344567_431;
   wire [7:0] v3_1645344567_432;
   wire [4:0] v3_1645344567_433;
   wire [7:0] v3_1645344567_434;
   wire [7:0] v3_1645344567_435;
   wire [7:0] v3_1645344567_436;
   wire [7:0] v3_1645344567_437;
   wire [7:0] v3_1645344567_438;
   wire [7:0] v3_1645344567_439;
   wire [7:0] v3_1645344567_440;
   wire [7:0] v3_1645344567_441;
   wire [7:0] v3_1645344567_442;
   wire [7:0] v3_1645344567_443;
   wire [7:0] v3_1645344567_444;
   wire [7:0] v3_1645344567_445;
   wire [7:0] v3_1645344567_446;
   wire [7:0] v3_1645344567_447;
   wire [7:0] v3_1645344567_448;
   wire [7:0] v3_1645344567_449;
   wire [7:0] v3_1645344567_450;
   wire v3_1645344567_451;

   // Output Net Declarations
   wire p;
   wire [2:0] coinOutNTD_50;
   wire [2:0] coinOutNTD_10;
   wire [2:0] coinOutNTD_5;
   wire [2:0] coinOutNTD_1;
   wire [1:0] itemTypeOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1645344567_0 = 1'b0; 
   assign v3_1645344567_23 = v3_1645344567_62 ? v3_1645344567_61 : v3_1645344567_24;
   assign v3_1645344567_24 = v3_1645344567_25;
   assign v3_1645344567_25 = v3_1645344567_60 ? v3_1645344567_56 : v3_1645344567_26;
   assign v3_1645344567_26 = v3_1645344567_55 ? v3_1645344567_54 : v3_1645344567_27;
   assign v3_1645344567_27 = v3_1645344567_53 ? v3_1645344567_32 : v3_1645344567_28;
   assign v3_1645344567_28 = v3_1645344567_51 ? v3_1645344567_43 : v3_1645344567_29;
   assign v3_1645344567_29 = v3_1645344567_41 ? v3_1645344567_32 : v3_1645344567_30;
   assign v3_1645344567_30 = v3_1645344567_39 ? v3_1645344567_32 : v3_1645344567_31;
   assign v3_1645344567_31 = v3_1645344567_37 ? v3_1645344567_33 : v3_1645344567_32;
   assign v3_1645344567_32 = v3_1645344567_8;
   assign v3_1645344567_33 = v3_1645344567_36 ? v3_1645344567_34 : v3_1645344567_32;
   assign v3_1645344567_34 = v3_1645344567_35;
   assign v3_1645344567_35 = 3'b000; 
   assign v3_1645344567_36 = v3_1645344567_21 == v3_1645344567_35;
   assign v3_1645344567_37 = v3_1645344567_18 >= v3_1645344567_38;
   assign v3_1645344567_38 = 8'b00000001; 
   assign v3_1645344567_39 = v3_1645344567_17 == v3_1645344567_40;
   assign v3_1645344567_40 = 2'b10; 
   assign v3_1645344567_41 = v3_1645344567_17 == v3_1645344567_42;
   assign v3_1645344567_42 = 2'b01; 
   assign v3_1645344567_43 = v3_1645344567_49 ? v3_1645344567_44 : v3_1645344567_32;
   assign v3_1645344567_44 = v3_1645344567_48 ? v3_1645344567_32 : v3_1645344567_45;
   assign v3_1645344567_45 = v3_1645344567_47;
   assign v3_1645344567_46 = 3'b001; 
   assign v3_1645344567_47 = v3_1645344567_8 + v3_1645344567_46;
   assign v3_1645344567_48 = v3_1645344567_19 == v3_1645344567_35;
   assign v3_1645344567_49 = v3_1645344567_18 >= v3_1645344567_50;
   assign v3_1645344567_50 = 8'b00110010; 
   assign v3_1645344567_51 = v3_1645344567_17 == v3_1645344567_52;
   assign v3_1645344567_52 = 2'b00; 
   assign v3_1645344567_53 = ~v3_1645344567_16;
   assign v3_1645344567_54 = v3_1645344567_35;
   assign v3_1645344567_55 = v3_1645344567_13 == v3_1645344567_52;
   assign v3_1645344567_56 = v3_1645344567_58 ? v3_1645344567_57 : v3_1645344567_32;
   assign v3_1645344567_57 = v3_1645344567_35;
   assign v3_1645344567_58 = ~v3_1645344567_59;
   assign v3_1645344567_59 = itemTypeIn == v3_1645344567_52;
   assign v3_1645344567_60 = v3_1645344567_13 == v3_1645344567_42;
   assign v3_1645344567_61 = v3_1645344567_35;
   assign v3_1645344567_62 = ~reset;
   assign v3_1645344567_63 = 3'b000; 
   assign v3_1645344567_64 = v3_1645344567_62 ? v3_1645344567_86 : v3_1645344567_65;
   assign v3_1645344567_65 = v3_1645344567_66;
   assign v3_1645344567_66 = v3_1645344567_60 ? v3_1645344567_84 : v3_1645344567_67;
   assign v3_1645344567_67 = v3_1645344567_55 ? v3_1645344567_83 : v3_1645344567_68;
   assign v3_1645344567_68 = v3_1645344567_53 ? v3_1645344567_73 : v3_1645344567_69;
   assign v3_1645344567_69 = v3_1645344567_51 ? v3_1645344567_73 : v3_1645344567_70;
   assign v3_1645344567_70 = v3_1645344567_41 ? v3_1645344567_76 : v3_1645344567_71;
   assign v3_1645344567_71 = v3_1645344567_39 ? v3_1645344567_73 : v3_1645344567_72;
   assign v3_1645344567_72 = v3_1645344567_37 ? v3_1645344567_74 : v3_1645344567_73;
   assign v3_1645344567_73 = v3_1645344567_9;
   assign v3_1645344567_74 = v3_1645344567_36 ? v3_1645344567_75 : v3_1645344567_73;
   assign v3_1645344567_75 = v3_1645344567_35;
   assign v3_1645344567_76 = v3_1645344567_81 ? v3_1645344567_77 : v3_1645344567_73;
   assign v3_1645344567_77 = v3_1645344567_80 ? v3_1645344567_73 : v3_1645344567_78;
   assign v3_1645344567_78 = v3_1645344567_79;
   assign v3_1645344567_79 = v3_1645344567_9 + v3_1645344567_46;
   assign v3_1645344567_80 = v3_1645344567_20 == v3_1645344567_35;
   assign v3_1645344567_81 = v3_1645344567_18 >= v3_1645344567_82;
   assign v3_1645344567_82 = 8'b00001010; 
   assign v3_1645344567_83 = v3_1645344567_35;
   assign v3_1645344567_84 = v3_1645344567_58 ? v3_1645344567_85 : v3_1645344567_73;
   assign v3_1645344567_85 = v3_1645344567_35;
   assign v3_1645344567_86 = v3_1645344567_35;
   assign v3_1645344567_87 = 3'b000; 
   assign v3_1645344567_88 = v3_1645344567_62 ? v3_1645344567_110 : v3_1645344567_89;
   assign v3_1645344567_89 = v3_1645344567_90;
   assign v3_1645344567_90 = v3_1645344567_60 ? v3_1645344567_108 : v3_1645344567_91;
   assign v3_1645344567_91 = v3_1645344567_55 ? v3_1645344567_107 : v3_1645344567_92;
   assign v3_1645344567_92 = v3_1645344567_53 ? v3_1645344567_97 : v3_1645344567_93;
   assign v3_1645344567_93 = v3_1645344567_51 ? v3_1645344567_97 : v3_1645344567_94;
   assign v3_1645344567_94 = v3_1645344567_41 ? v3_1645344567_97 : v3_1645344567_95;
   assign v3_1645344567_95 = v3_1645344567_39 ? v3_1645344567_100 : v3_1645344567_96;
   assign v3_1645344567_96 = v3_1645344567_37 ? v3_1645344567_98 : v3_1645344567_97;
   assign v3_1645344567_97 = v3_1645344567_10;
   assign v3_1645344567_98 = v3_1645344567_36 ? v3_1645344567_99 : v3_1645344567_97;
   assign v3_1645344567_99 = v3_1645344567_35;
   assign v3_1645344567_100 = v3_1645344567_105 ? v3_1645344567_101 : v3_1645344567_97;
   assign v3_1645344567_101 = v3_1645344567_104 ? v3_1645344567_97 : v3_1645344567_102;
   assign v3_1645344567_102 = v3_1645344567_103;
   assign v3_1645344567_103 = v3_1645344567_10 + v3_1645344567_46;
   assign v3_1645344567_104 = v3_1645344567_22 == v3_1645344567_35;
   assign v3_1645344567_105 = v3_1645344567_18 >= v3_1645344567_106;
   assign v3_1645344567_106 = 8'b00000101; 
   assign v3_1645344567_107 = v3_1645344567_35;
   assign v3_1645344567_108 = v3_1645344567_58 ? v3_1645344567_109 : v3_1645344567_97;
   assign v3_1645344567_109 = v3_1645344567_35;
   assign v3_1645344567_110 = v3_1645344567_35;
   assign v3_1645344567_111 = 3'b000; 
   assign v3_1645344567_112 = v3_1645344567_62 ? v3_1645344567_129 : v3_1645344567_113;
   assign v3_1645344567_113 = v3_1645344567_114;
   assign v3_1645344567_114 = v3_1645344567_60 ? v3_1645344567_127 : v3_1645344567_115;
   assign v3_1645344567_115 = v3_1645344567_55 ? v3_1645344567_126 : v3_1645344567_116;
   assign v3_1645344567_116 = v3_1645344567_53 ? v3_1645344567_121 : v3_1645344567_117;
   assign v3_1645344567_117 = v3_1645344567_51 ? v3_1645344567_121 : v3_1645344567_118;
   assign v3_1645344567_118 = v3_1645344567_41 ? v3_1645344567_121 : v3_1645344567_119;
   assign v3_1645344567_119 = v3_1645344567_39 ? v3_1645344567_121 : v3_1645344567_120;
   assign v3_1645344567_120 = v3_1645344567_37 ? v3_1645344567_122 : v3_1645344567_121;
   assign v3_1645344567_121 = v3_1645344567_11;
   assign v3_1645344567_122 = v3_1645344567_36 ? v3_1645344567_125 : v3_1645344567_123;
   assign v3_1645344567_123 = v3_1645344567_124;
   assign v3_1645344567_124 = v3_1645344567_11 + v3_1645344567_46;
   assign v3_1645344567_125 = v3_1645344567_35;
   assign v3_1645344567_126 = v3_1645344567_35;
   assign v3_1645344567_127 = v3_1645344567_58 ? v3_1645344567_128 : v3_1645344567_121;
   assign v3_1645344567_128 = v3_1645344567_35;
   assign v3_1645344567_129 = v3_1645344567_35;
   assign v3_1645344567_130 = 3'b000; 
   assign v3_1645344567_131 = v3_1645344567_62 ? v3_1645344567_150 : v3_1645344567_132;
   assign v3_1645344567_132 = v3_1645344567_133;
   assign v3_1645344567_133 = v3_1645344567_60 ? v3_1645344567_148 : v3_1645344567_134;
   assign v3_1645344567_134 = v3_1645344567_55 ? v3_1645344567_147 : v3_1645344567_135;
   assign v3_1645344567_135 = v3_1645344567_53 ? v3_1645344567_143 : v3_1645344567_136;
   assign v3_1645344567_136 = v3_1645344567_51 ? v3_1645344567_140 : v3_1645344567_137;
   assign v3_1645344567_137 = v3_1645344567_41 ? v3_1645344567_140 : v3_1645344567_138;
   assign v3_1645344567_138 = v3_1645344567_39 ? v3_1645344567_140 : v3_1645344567_139;
   assign v3_1645344567_139 = v3_1645344567_37 ? v3_1645344567_141 : v3_1645344567_140;
   assign v3_1645344567_140 = v3_1645344567_12;
   assign v3_1645344567_141 = v3_1645344567_36 ? v3_1645344567_142 : v3_1645344567_140;
   assign v3_1645344567_142 = v3_1645344567_52;
   assign v3_1645344567_143 = v3_1645344567_145 ? v3_1645344567_144 : v3_1645344567_140;
   assign v3_1645344567_144 = v3_1645344567_52;
   assign v3_1645344567_145 = ~v3_1645344567_146;
   assign v3_1645344567_146 = v3_1645344567_15 >= v3_1645344567_18;
   assign v3_1645344567_147 = v3_1645344567_52;
   assign v3_1645344567_148 = v3_1645344567_58 ? v3_1645344567_149 : v3_1645344567_140;
   assign v3_1645344567_149 = itemTypeIn;
   assign v3_1645344567_150 = v3_1645344567_52;
   assign v3_1645344567_151 = 2'b00; 
   assign v3_1645344567_152 = v3_1645344567_62 ? v3_1645344567_168 : v3_1645344567_153;
   assign v3_1645344567_153 = v3_1645344567_154;
   assign v3_1645344567_154 = v3_1645344567_60 ? v3_1645344567_166 : v3_1645344567_155;
   assign v3_1645344567_155 = v3_1645344567_55 ? v3_1645344567_165 : v3_1645344567_156;
   assign v3_1645344567_156 = v3_1645344567_53 ? v3_1645344567_163 : v3_1645344567_157;
   assign v3_1645344567_157 = v3_1645344567_51 ? v3_1645344567_163 : v3_1645344567_158;
   assign v3_1645344567_158 = v3_1645344567_41 ? v3_1645344567_163 : v3_1645344567_159;
   assign v3_1645344567_159 = v3_1645344567_39 ? v3_1645344567_163 : v3_1645344567_160;
   assign v3_1645344567_160 = v3_1645344567_37 ? v3_1645344567_162 : v3_1645344567_161;
   assign v3_1645344567_161 = v3_1645344567_52;
   assign v3_1645344567_162 = v3_1645344567_36 ? v3_1645344567_164 : v3_1645344567_163;
   assign v3_1645344567_163 = v3_1645344567_13;
   assign v3_1645344567_164 = v3_1645344567_52;
   assign v3_1645344567_165 = v3_1645344567_42;
   assign v3_1645344567_166 = v3_1645344567_58 ? v3_1645344567_167 : v3_1645344567_163;
   assign v3_1645344567_167 = v3_1645344567_40;
   assign v3_1645344567_168 = v3_1645344567_42;
   assign v3_1645344567_169 = 2'b00; 
   assign v3_1645344567_170 = v3_1645344567_62 ? v3_1645344567_172 : v3_1645344567_171;
   assign v3_1645344567_171 = v3_1645344567_14;
   assign v3_1645344567_172 = v3_1645344567_173;
   assign v3_1645344567_173 = 1'b1; 
   assign v3_1645344567_174 = 1'b0; 
   assign v3_1645344567_175 = v3_1645344567_62 ? v3_1645344567_203 : v3_1645344567_176;
   assign v3_1645344567_176 = v3_1645344567_177;
   assign v3_1645344567_177 = v3_1645344567_60 ? v3_1645344567_179 : v3_1645344567_178;
   assign v3_1645344567_178 = v3_1645344567_15;
   assign v3_1645344567_179 = v3_1645344567_58 ? v3_1645344567_180 : v3_1645344567_178;
   assign v3_1645344567_180 = v3_1645344567_202;
   assign v3_1645344567_181 = v3_1645344567_197;
   assign v3_1645344567_182 = v3_1645344567_192;
   assign v3_1645344567_183 = v3_1645344567_187;
   assign v3_1645344567_184 = v3_1645344567_186;
   assign v3_1645344567_185 = 6'b000000; 
   assign v3_1645344567_186 = {v3_1645344567_185, coinInNTD_50};
   assign v3_1645344567_187 = v3_1645344567_50 * v3_1645344567_184;
   assign v3_1645344567_188 = v3_1645344567_191;
   assign v3_1645344567_189 = v3_1645344567_190;
   assign v3_1645344567_190 = {v3_1645344567_185, coinInNTD_10};
   assign v3_1645344567_191 = v3_1645344567_82 * v3_1645344567_189;
   assign v3_1645344567_192 = v3_1645344567_183 + v3_1645344567_188;
   assign v3_1645344567_193 = v3_1645344567_196;
   assign v3_1645344567_194 = v3_1645344567_195;
   assign v3_1645344567_195 = {v3_1645344567_185, coinInNTD_5};
   assign v3_1645344567_196 = v3_1645344567_106 * v3_1645344567_194;
   assign v3_1645344567_197 = v3_1645344567_182 + v3_1645344567_193;
   assign v3_1645344567_198 = v3_1645344567_201;
   assign v3_1645344567_199 = v3_1645344567_200;
   assign v3_1645344567_200 = {v3_1645344567_185, coinInNTD_1};
   assign v3_1645344567_201 = v3_1645344567_38 * v3_1645344567_199;
   assign v3_1645344567_202 = v3_1645344567_181 + v3_1645344567_198;
   assign v3_1645344567_203 = v3_1645344567_204;
   assign v3_1645344567_204 = 8'b00000000; 
   assign v3_1645344567_205 = 8'b00000000; 
   assign v3_1645344567_206 = v3_1645344567_62 ? v3_1645344567_218 : v3_1645344567_207;
   assign v3_1645344567_207 = v3_1645344567_208;
   assign v3_1645344567_208 = v3_1645344567_60 ? v3_1645344567_215 : v3_1645344567_209;
   assign v3_1645344567_209 = v3_1645344567_55 ? v3_1645344567_211 : v3_1645344567_210;
   assign v3_1645344567_210 = v3_1645344567_53 ? v3_1645344567_212 : v3_1645344567_211;
   assign v3_1645344567_211 = v3_1645344567_16;
   assign v3_1645344567_212 = v3_1645344567_145 ? v3_1645344567_214 : v3_1645344567_213;
   assign v3_1645344567_213 = v3_1645344567_173;
   assign v3_1645344567_214 = v3_1645344567_173;
   assign v3_1645344567_215 = v3_1645344567_58 ? v3_1645344567_216 : v3_1645344567_211;
   assign v3_1645344567_216 = v3_1645344567_217;
   assign v3_1645344567_217 = 1'b0; 
   assign v3_1645344567_218 = v3_1645344567_217;
   assign v3_1645344567_219 = 1'b0; 
   assign v3_1645344567_220 = v3_1645344567_62 ? v3_1645344567_247 : v3_1645344567_221;
   assign v3_1645344567_221 = v3_1645344567_222;
   assign v3_1645344567_222 = v3_1645344567_60 ? v3_1645344567_245 : v3_1645344567_223;
   assign v3_1645344567_223 = v3_1645344567_55 ? v3_1645344567_229 : v3_1645344567_224;
   assign v3_1645344567_224 = v3_1645344567_53 ? v3_1645344567_229 : v3_1645344567_225;
   assign v3_1645344567_225 = v3_1645344567_51 ? v3_1645344567_241 : v3_1645344567_226;
   assign v3_1645344567_226 = v3_1645344567_41 ? v3_1645344567_237 : v3_1645344567_227;
   assign v3_1645344567_227 = v3_1645344567_39 ? v3_1645344567_232 : v3_1645344567_228;
   assign v3_1645344567_228 = v3_1645344567_37 ? v3_1645344567_230 : v3_1645344567_229;
   assign v3_1645344567_229 = v3_1645344567_17;
   assign v3_1645344567_230 = v3_1645344567_36 ? v3_1645344567_231 : v3_1645344567_229;
   assign v3_1645344567_231 = v3_1645344567_52;
   assign v3_1645344567_232 = v3_1645344567_105 ? v3_1645344567_235 : v3_1645344567_233;
   assign v3_1645344567_233 = v3_1645344567_234;
   assign v3_1645344567_234 = 2'b11; 
   assign v3_1645344567_235 = v3_1645344567_104 ? v3_1645344567_236 : v3_1645344567_229;
   assign v3_1645344567_236 = v3_1645344567_234;
   assign v3_1645344567_237 = v3_1645344567_81 ? v3_1645344567_239 : v3_1645344567_238;
   assign v3_1645344567_238 = v3_1645344567_40;
   assign v3_1645344567_239 = v3_1645344567_80 ? v3_1645344567_240 : v3_1645344567_229;
   assign v3_1645344567_240 = v3_1645344567_40;
   assign v3_1645344567_241 = v3_1645344567_49 ? v3_1645344567_243 : v3_1645344567_242;
   assign v3_1645344567_242 = v3_1645344567_42;
   assign v3_1645344567_243 = v3_1645344567_48 ? v3_1645344567_244 : v3_1645344567_229;
   assign v3_1645344567_244 = v3_1645344567_42;
   assign v3_1645344567_245 = v3_1645344567_58 ? v3_1645344567_246 : v3_1645344567_229;
   assign v3_1645344567_246 = v3_1645344567_52;
   assign v3_1645344567_247 = v3_1645344567_52;
   assign v3_1645344567_248 = 2'b00; 
   assign v3_1645344567_249 = v3_1645344567_62 ? v3_1645344567_289 : v3_1645344567_250;
   assign v3_1645344567_250 = v3_1645344567_251;
   assign v3_1645344567_251 = v3_1645344567_60 ? v3_1645344567_279 : v3_1645344567_252;
   assign v3_1645344567_252 = v3_1645344567_55 ? v3_1645344567_258 : v3_1645344567_253;
   assign v3_1645344567_253 = v3_1645344567_53 ? v3_1645344567_275 : v3_1645344567_254;
   assign v3_1645344567_254 = v3_1645344567_51 ? v3_1645344567_271 : v3_1645344567_255;
   assign v3_1645344567_255 = v3_1645344567_41 ? v3_1645344567_267 : v3_1645344567_256;
   assign v3_1645344567_256 = v3_1645344567_39 ? v3_1645344567_263 : v3_1645344567_257;
   assign v3_1645344567_257 = v3_1645344567_37 ? v3_1645344567_259 : v3_1645344567_258;
   assign v3_1645344567_258 = v3_1645344567_18;
   assign v3_1645344567_259 = v3_1645344567_36 ? v3_1645344567_262 : v3_1645344567_260;
   assign v3_1645344567_260 = v3_1645344567_261;
   assign v3_1645344567_261 = v3_1645344567_18 - v3_1645344567_38;
   assign v3_1645344567_262 = v3_1645344567_15;
   assign v3_1645344567_263 = v3_1645344567_105 ? v3_1645344567_264 : v3_1645344567_258;
   assign v3_1645344567_264 = v3_1645344567_104 ? v3_1645344567_258 : v3_1645344567_265;
   assign v3_1645344567_265 = v3_1645344567_266;
   assign v3_1645344567_266 = v3_1645344567_18 - v3_1645344567_106;
   assign v3_1645344567_267 = v3_1645344567_81 ? v3_1645344567_268 : v3_1645344567_258;
   assign v3_1645344567_268 = v3_1645344567_80 ? v3_1645344567_258 : v3_1645344567_269;
   assign v3_1645344567_269 = v3_1645344567_270;
   assign v3_1645344567_270 = v3_1645344567_18 - v3_1645344567_82;
   assign v3_1645344567_271 = v3_1645344567_49 ? v3_1645344567_272 : v3_1645344567_258;
   assign v3_1645344567_272 = v3_1645344567_48 ? v3_1645344567_258 : v3_1645344567_273;
   assign v3_1645344567_273 = v3_1645344567_274;
   assign v3_1645344567_274 = v3_1645344567_18 - v3_1645344567_50;
   assign v3_1645344567_275 = v3_1645344567_145 ? v3_1645344567_278 : v3_1645344567_276;
   assign v3_1645344567_276 = v3_1645344567_277;
   assign v3_1645344567_277 = v3_1645344567_15 - v3_1645344567_18;
   assign v3_1645344567_278 = v3_1645344567_15;
   assign v3_1645344567_279 = v3_1645344567_58 ? v3_1645344567_280 : v3_1645344567_258;
   assign v3_1645344567_280 = v3_1645344567_288 ? v3_1645344567_287 : v3_1645344567_281;
   assign v3_1645344567_281 = v3_1645344567_286 ? v3_1645344567_285 : v3_1645344567_282;
   assign v3_1645344567_282 = v3_1645344567_284 ? v3_1645344567_283 : v3_1645344567_204;
   assign v3_1645344567_283 = 8'b00010110; 
   assign v3_1645344567_284 = itemTypeIn == v3_1645344567_234;
   assign v3_1645344567_285 = 8'b00001111; 
   assign v3_1645344567_286 = itemTypeIn == v3_1645344567_40;
   assign v3_1645344567_287 = 8'b00001000; 
   assign v3_1645344567_288 = itemTypeIn == v3_1645344567_42;
   assign v3_1645344567_289 = v3_1645344567_204;
   assign v3_1645344567_290 = 8'b00000000; 
   assign v3_1645344567_291 = v3_1645344567_62 ? v3_1645344567_323 : v3_1645344567_292;
   assign v3_1645344567_292 = v3_1645344567_293;
   assign v3_1645344567_293 = v3_1645344567_60 ? v3_1645344567_308 : v3_1645344567_294;
   assign v3_1645344567_294 = v3_1645344567_55 ? v3_1645344567_300 : v3_1645344567_295;
   assign v3_1645344567_295 = v3_1645344567_53 ? v3_1645344567_300 : v3_1645344567_296;
   assign v3_1645344567_296 = v3_1645344567_51 ? v3_1645344567_304 : v3_1645344567_297;
   assign v3_1645344567_297 = v3_1645344567_41 ? v3_1645344567_300 : v3_1645344567_298;
   assign v3_1645344567_298 = v3_1645344567_39 ? v3_1645344567_300 : v3_1645344567_299;
   assign v3_1645344567_299 = v3_1645344567_37 ? v3_1645344567_301 : v3_1645344567_300;
   assign v3_1645344567_300 = v3_1645344567_19;
   assign v3_1645344567_301 = v3_1645344567_36 ? v3_1645344567_302 : v3_1645344567_300;
   assign v3_1645344567_302 = v3_1645344567_303;
   assign v3_1645344567_303 = v3_1645344567_19 + v3_1645344567_8;
   assign v3_1645344567_304 = v3_1645344567_49 ? v3_1645344567_305 : v3_1645344567_300;
   assign v3_1645344567_305 = v3_1645344567_48 ? v3_1645344567_300 : v3_1645344567_306;
   assign v3_1645344567_306 = v3_1645344567_307;
   assign v3_1645344567_307 = v3_1645344567_19 - v3_1645344567_46;
   assign v3_1645344567_308 = v3_1645344567_58 ? v3_1645344567_309 : v3_1645344567_300;
   assign v3_1645344567_309 = v3_1645344567_315 ? v3_1645344567_314 : v3_1645344567_310;
   assign v3_1645344567_310 = v3_1645344567_313;
   assign v3_1645344567_311 = v3_1645344567_312;
   assign v3_1645344567_312 = {v3_1645344567_217, coinInNTD_50};
   assign v3_1645344567_313 = v3_1645344567_19 + v3_1645344567_311;
   assign v3_1645344567_314 = 3'b111; 
   assign v3_1645344567_315 = v3_1645344567_316 >= v3_1645344567_322;
   assign v3_1645344567_316 = v3_1645344567_321;
   assign v3_1645344567_317 = v3_1645344567_318;
   assign v3_1645344567_318 = {v3_1645344567_217, v3_1645344567_19};
   assign v3_1645344567_319 = v3_1645344567_320;
   assign v3_1645344567_320 = {v3_1645344567_52, coinInNTD_50};
   assign v3_1645344567_321 = v3_1645344567_317 + v3_1645344567_319;
   assign v3_1645344567_322 = 4'b0111; 
   assign v3_1645344567_323 = v3_1645344567_324;
   assign v3_1645344567_324 = 3'b010; 
   assign v3_1645344567_325 = 3'b000; 
   assign v3_1645344567_326 = v3_1645344567_62 ? v3_1645344567_356 : v3_1645344567_327;
   assign v3_1645344567_327 = v3_1645344567_328;
   assign v3_1645344567_328 = v3_1645344567_60 ? v3_1645344567_343 : v3_1645344567_329;
   assign v3_1645344567_329 = v3_1645344567_55 ? v3_1645344567_335 : v3_1645344567_330;
   assign v3_1645344567_330 = v3_1645344567_53 ? v3_1645344567_335 : v3_1645344567_331;
   assign v3_1645344567_331 = v3_1645344567_51 ? v3_1645344567_335 : v3_1645344567_332;
   assign v3_1645344567_332 = v3_1645344567_41 ? v3_1645344567_339 : v3_1645344567_333;
   assign v3_1645344567_333 = v3_1645344567_39 ? v3_1645344567_335 : v3_1645344567_334;
   assign v3_1645344567_334 = v3_1645344567_37 ? v3_1645344567_336 : v3_1645344567_335;
   assign v3_1645344567_335 = v3_1645344567_20;
   assign v3_1645344567_336 = v3_1645344567_36 ? v3_1645344567_337 : v3_1645344567_335;
   assign v3_1645344567_337 = v3_1645344567_338;
   assign v3_1645344567_338 = v3_1645344567_20 + v3_1645344567_9;
   assign v3_1645344567_339 = v3_1645344567_81 ? v3_1645344567_340 : v3_1645344567_335;
   assign v3_1645344567_340 = v3_1645344567_80 ? v3_1645344567_335 : v3_1645344567_341;
   assign v3_1645344567_341 = v3_1645344567_342;
   assign v3_1645344567_342 = v3_1645344567_20 - v3_1645344567_46;
   assign v3_1645344567_343 = v3_1645344567_58 ? v3_1645344567_344 : v3_1645344567_335;
   assign v3_1645344567_344 = v3_1645344567_349 ? v3_1645344567_314 : v3_1645344567_345;
   assign v3_1645344567_345 = v3_1645344567_348;
   assign v3_1645344567_346 = v3_1645344567_347;
   assign v3_1645344567_347 = {v3_1645344567_217, coinInNTD_10};
   assign v3_1645344567_348 = v3_1645344567_20 + v3_1645344567_346;
   assign v3_1645344567_349 = v3_1645344567_350 >= v3_1645344567_322;
   assign v3_1645344567_350 = v3_1645344567_355;
   assign v3_1645344567_351 = v3_1645344567_352;
   assign v3_1645344567_352 = {v3_1645344567_217, v3_1645344567_20};
   assign v3_1645344567_353 = v3_1645344567_354;
   assign v3_1645344567_354 = {v3_1645344567_52, coinInNTD_10};
   assign v3_1645344567_355 = v3_1645344567_351 + v3_1645344567_353;
   assign v3_1645344567_356 = v3_1645344567_324;
   assign v3_1645344567_357 = 3'b000; 
   assign v3_1645344567_358 = v3_1645344567_62 ? v3_1645344567_386 : v3_1645344567_359;
   assign v3_1645344567_359 = v3_1645344567_360;
   assign v3_1645344567_360 = v3_1645344567_60 ? v3_1645344567_373 : v3_1645344567_361;
   assign v3_1645344567_361 = v3_1645344567_55 ? v3_1645344567_367 : v3_1645344567_362;
   assign v3_1645344567_362 = v3_1645344567_53 ? v3_1645344567_367 : v3_1645344567_363;
   assign v3_1645344567_363 = v3_1645344567_51 ? v3_1645344567_367 : v3_1645344567_364;
   assign v3_1645344567_364 = v3_1645344567_41 ? v3_1645344567_367 : v3_1645344567_365;
   assign v3_1645344567_365 = v3_1645344567_39 ? v3_1645344567_367 : v3_1645344567_366;
   assign v3_1645344567_366 = v3_1645344567_37 ? v3_1645344567_368 : v3_1645344567_367;
   assign v3_1645344567_367 = v3_1645344567_21;
   assign v3_1645344567_368 = v3_1645344567_36 ? v3_1645344567_371 : v3_1645344567_369;
   assign v3_1645344567_369 = v3_1645344567_370;
   assign v3_1645344567_370 = v3_1645344567_21 - v3_1645344567_46;
   assign v3_1645344567_371 = v3_1645344567_372;
   assign v3_1645344567_372 = v3_1645344567_21 + v3_1645344567_11;
   assign v3_1645344567_373 = v3_1645344567_58 ? v3_1645344567_374 : v3_1645344567_367;
   assign v3_1645344567_374 = v3_1645344567_379 ? v3_1645344567_314 : v3_1645344567_375;
   assign v3_1645344567_375 = v3_1645344567_378;
   assign v3_1645344567_376 = v3_1645344567_377;
   assign v3_1645344567_377 = {v3_1645344567_217, coinInNTD_1};
   assign v3_1645344567_378 = v3_1645344567_21 + v3_1645344567_376;
   assign v3_1645344567_379 = v3_1645344567_380 >= v3_1645344567_322;
   assign v3_1645344567_380 = v3_1645344567_385;
   assign v3_1645344567_381 = v3_1645344567_382;
   assign v3_1645344567_382 = {v3_1645344567_217, v3_1645344567_21};
   assign v3_1645344567_383 = v3_1645344567_384;
   assign v3_1645344567_384 = {v3_1645344567_52, coinInNTD_1};
   assign v3_1645344567_385 = v3_1645344567_381 + v3_1645344567_383;
   assign v3_1645344567_386 = v3_1645344567_324;
   assign v3_1645344567_387 = 3'b000; 
   assign v3_1645344567_388 = v3_1645344567_62 ? v3_1645344567_418 : v3_1645344567_389;
   assign v3_1645344567_389 = v3_1645344567_390;
   assign v3_1645344567_390 = v3_1645344567_60 ? v3_1645344567_405 : v3_1645344567_391;
   assign v3_1645344567_391 = v3_1645344567_55 ? v3_1645344567_397 : v3_1645344567_392;
   assign v3_1645344567_392 = v3_1645344567_53 ? v3_1645344567_397 : v3_1645344567_393;
   assign v3_1645344567_393 = v3_1645344567_51 ? v3_1645344567_397 : v3_1645344567_394;
   assign v3_1645344567_394 = v3_1645344567_41 ? v3_1645344567_397 : v3_1645344567_395;
   assign v3_1645344567_395 = v3_1645344567_39 ? v3_1645344567_401 : v3_1645344567_396;
   assign v3_1645344567_396 = v3_1645344567_37 ? v3_1645344567_398 : v3_1645344567_397;
   assign v3_1645344567_397 = v3_1645344567_22;
   assign v3_1645344567_398 = v3_1645344567_36 ? v3_1645344567_399 : v3_1645344567_397;
   assign v3_1645344567_399 = v3_1645344567_400;
   assign v3_1645344567_400 = v3_1645344567_22 + v3_1645344567_10;
   assign v3_1645344567_401 = v3_1645344567_105 ? v3_1645344567_402 : v3_1645344567_397;
   assign v3_1645344567_402 = v3_1645344567_104 ? v3_1645344567_397 : v3_1645344567_403;
   assign v3_1645344567_403 = v3_1645344567_404;
   assign v3_1645344567_404 = v3_1645344567_22 - v3_1645344567_46;
   assign v3_1645344567_405 = v3_1645344567_58 ? v3_1645344567_406 : v3_1645344567_397;
   assign v3_1645344567_406 = v3_1645344567_411 ? v3_1645344567_314 : v3_1645344567_407;
   assign v3_1645344567_407 = v3_1645344567_410;
   assign v3_1645344567_408 = v3_1645344567_409;
   assign v3_1645344567_409 = {v3_1645344567_217, coinInNTD_5};
   assign v3_1645344567_410 = v3_1645344567_22 + v3_1645344567_408;
   assign v3_1645344567_411 = v3_1645344567_412 >= v3_1645344567_322;
   assign v3_1645344567_412 = v3_1645344567_417;
   assign v3_1645344567_413 = v3_1645344567_414;
   assign v3_1645344567_414 = {v3_1645344567_217, v3_1645344567_22};
   assign v3_1645344567_415 = v3_1645344567_416;
   assign v3_1645344567_416 = {v3_1645344567_52, coinInNTD_5};
   assign v3_1645344567_417 = v3_1645344567_413 + v3_1645344567_415;
   assign v3_1645344567_418 = v3_1645344567_324;
   assign v3_1645344567_419 = 3'b000; 
   assign v3_1645344567_420 = v3_1645344567_451;
   assign v3_1645344567_421 = v3_1645344567_425;
   assign v3_1645344567_422 = v3_1645344567_423;
   assign v3_1645344567_423 = v3_1645344567_14 & v3_1645344567_55;
   assign v3_1645344567_424 = v3_1645344567_12 == v3_1645344567_52;
   assign v3_1645344567_425 = v3_1645344567_422 & v3_1645344567_424;
   assign v3_1645344567_426 = ~v3_1645344567_427;
   assign v3_1645344567_427 = v3_1645344567_428 == v3_1645344567_15;
   assign v3_1645344567_428 = v3_1645344567_450;
   assign v3_1645344567_429 = v3_1645344567_445;
   assign v3_1645344567_430 = v3_1645344567_440;
   assign v3_1645344567_431 = v3_1645344567_435;
   assign v3_1645344567_432 = v3_1645344567_434;
   assign v3_1645344567_433 = 5'b00000; 
   assign v3_1645344567_434 = {v3_1645344567_433, v3_1645344567_8};
   assign v3_1645344567_435 = v3_1645344567_50 * v3_1645344567_432;
   assign v3_1645344567_436 = v3_1645344567_439;
   assign v3_1645344567_437 = v3_1645344567_438;
   assign v3_1645344567_438 = {v3_1645344567_433, v3_1645344567_9};
   assign v3_1645344567_439 = v3_1645344567_82 * v3_1645344567_437;
   assign v3_1645344567_440 = v3_1645344567_431 + v3_1645344567_436;
   assign v3_1645344567_441 = v3_1645344567_444;
   assign v3_1645344567_442 = v3_1645344567_443;
   assign v3_1645344567_443 = {v3_1645344567_433, v3_1645344567_10};
   assign v3_1645344567_444 = v3_1645344567_106 * v3_1645344567_442;
   assign v3_1645344567_445 = v3_1645344567_430 + v3_1645344567_441;
   assign v3_1645344567_446 = v3_1645344567_449;
   assign v3_1645344567_447 = v3_1645344567_448;
   assign v3_1645344567_448 = {v3_1645344567_433, v3_1645344567_11};
   assign v3_1645344567_449 = v3_1645344567_38 * v3_1645344567_447;
   assign v3_1645344567_450 = v3_1645344567_429 + v3_1645344567_446;
   assign v3_1645344567_451 = v3_1645344567_421 & v3_1645344567_426;

   // Output Net Assignments
   assign p = v3_1645344567_420;
   assign coinOutNTD_50 = v3_1645344567_8;
   assign coinOutNTD_10 = v3_1645344567_9;
   assign coinOutNTD_5 = v3_1645344567_10;
   assign coinOutNTD_1 = v3_1645344567_11;
   assign itemTypeOut = v3_1645344567_12;
   assign serviceTypeOut = v3_1645344567_13;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1645344567_8 <= v3_1645344567_23;
      v3_1645344567_9 <= v3_1645344567_64;
      v3_1645344567_10 <= v3_1645344567_88;
      v3_1645344567_11 <= v3_1645344567_112;
      v3_1645344567_12 <= v3_1645344567_131;
      v3_1645344567_13 <= v3_1645344567_152;
      v3_1645344567_14 <= v3_1645344567_170;
      v3_1645344567_15 <= v3_1645344567_175;
      v3_1645344567_16 <= v3_1645344567_206;
      v3_1645344567_17 <= v3_1645344567_220;
      v3_1645344567_18 <= v3_1645344567_249;
      v3_1645344567_19 <= v3_1645344567_291;
      v3_1645344567_20 <= v3_1645344567_326;
      v3_1645344567_21 <= v3_1645344567_358;
      v3_1645344567_22 <= v3_1645344567_388;
   end
endmodule
