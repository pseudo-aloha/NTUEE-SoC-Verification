// RTL (Verilog) generated @ Mon Mar  7 14:51:29 2022 by V3 
//               compiled @ Feb 20 2022 16:07:45
// Internal nets are renamed with prefix "v3_1646635889_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire id0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] coinOutNTD_50;
   reg [2:0] coinOutNTD_10;
   reg [2:0] coinOutNTD_5;
   reg [2:0] coinOutNTD_1;
   reg [1:0] itemTypeOut;
   reg [1:0] serviceTypeOut;
   reg initialized;
   reg [7:0] inputValue;
   reg exchangeReady;
   reg [1:0] serviceCoinType;
   reg [7:0] serviceValue;
   reg [2:0] countNTD_50;
   reg [2:0] countNTD_10;
   reg [2:0] countNTD_1;
   reg [2:0] countNTD_5;
   wire [2:0] v3_1646635889_23;
   wire [2:0] v3_1646635889_24;
   wire [2:0] coinOutNTD_50_w;
   wire [2:0] v3_1646635889_26;
   wire [2:0] v3_1646635889_27;
   wire [2:0] v3_1646635889_28;
   wire [2:0] v3_1646635889_29;
   wire [2:0] v3_1646635889_30;
   wire [2:0] v3_1646635889_31;
   wire [2:0] v3_1646635889_32;
   wire [2:0] v3_1646635889_33;
   wire [2:0] v3_1646635889_34;
   wire [2:0] v3_1646635889_35;
   wire v3_1646635889_36;
   wire v3_1646635889_37;
   wire [7:0] v3_1646635889_38;
   wire v3_1646635889_39;
   wire [1:0] v3_1646635889_40;
   wire v3_1646635889_41;
   wire [1:0] v3_1646635889_42;
   wire [2:0] v3_1646635889_43;
   wire [2:0] v3_1646635889_44;
   wire [2:0] v3_1646635889_45;
   wire [2:0] v3_1646635889_46;
   wire [2:0] v3_1646635889_47;
   wire v3_1646635889_48;
   wire v3_1646635889_49;
   wire [7:0] v3_1646635889_50;
   wire v3_1646635889_51;
   wire [1:0] v3_1646635889_52;
   wire v3_1646635889_53;
   wire [2:0] v3_1646635889_54;
   wire v3_1646635889_55;
   wire [2:0] v3_1646635889_56;
   wire [2:0] v3_1646635889_57;
   wire v3_1646635889_58;
   wire v3_1646635889_59;
   wire v3_1646635889_60;
   wire [2:0] v3_1646635889_61;
   wire v3_1646635889_62;
   wire [2:0] v3_1646635889_63;
   wire [2:0] v3_1646635889_64;
   wire [2:0] v3_1646635889_65;
   wire [2:0] coinOutNTD_10_w;
   wire [2:0] v3_1646635889_67;
   wire [2:0] v3_1646635889_68;
   wire [2:0] v3_1646635889_69;
   wire [2:0] v3_1646635889_70;
   wire [2:0] v3_1646635889_71;
   wire [2:0] v3_1646635889_72;
   wire [2:0] v3_1646635889_73;
   wire [2:0] v3_1646635889_74;
   wire [2:0] v3_1646635889_75;
   wire [2:0] v3_1646635889_76;
   wire [2:0] v3_1646635889_77;
   wire [2:0] v3_1646635889_78;
   wire [2:0] v3_1646635889_79;
   wire v3_1646635889_80;
   wire v3_1646635889_81;
   wire [7:0] v3_1646635889_82;
   wire [2:0] v3_1646635889_83;
   wire [2:0] v3_1646635889_84;
   wire [2:0] v3_1646635889_85;
   wire [2:0] v3_1646635889_86;
   wire [2:0] v3_1646635889_87;
   wire [2:0] v3_1646635889_88;
   wire [2:0] v3_1646635889_89;
   wire [2:0] coinOutNTD_5_w;
   wire [2:0] v3_1646635889_91;
   wire [2:0] v3_1646635889_92;
   wire [2:0] v3_1646635889_93;
   wire [2:0] v3_1646635889_94;
   wire [2:0] v3_1646635889_95;
   wire [2:0] v3_1646635889_96;
   wire [2:0] v3_1646635889_97;
   wire [2:0] v3_1646635889_98;
   wire [2:0] v3_1646635889_99;
   wire [2:0] v3_1646635889_100;
   wire [2:0] v3_1646635889_101;
   wire [2:0] v3_1646635889_102;
   wire [2:0] v3_1646635889_103;
   wire v3_1646635889_104;
   wire v3_1646635889_105;
   wire [7:0] v3_1646635889_106;
   wire [2:0] v3_1646635889_107;
   wire [2:0] v3_1646635889_108;
   wire [2:0] v3_1646635889_109;
   wire [2:0] v3_1646635889_110;
   wire [2:0] v3_1646635889_111;
   wire [2:0] v3_1646635889_112;
   wire [2:0] v3_1646635889_113;
   wire [2:0] coinOutNTD_1_w;
   wire [2:0] v3_1646635889_115;
   wire [2:0] v3_1646635889_116;
   wire [2:0] v3_1646635889_117;
   wire [2:0] v3_1646635889_118;
   wire [2:0] v3_1646635889_119;
   wire [2:0] v3_1646635889_120;
   wire [2:0] v3_1646635889_121;
   wire [2:0] v3_1646635889_122;
   wire [2:0] v3_1646635889_123;
   wire [2:0] v3_1646635889_124;
   wire [2:0] v3_1646635889_125;
   wire [2:0] v3_1646635889_126;
   wire [2:0] v3_1646635889_127;
   wire [2:0] v3_1646635889_128;
   wire [2:0] v3_1646635889_129;
   wire [2:0] v3_1646635889_130;
   wire [1:0] v3_1646635889_131;
   wire [1:0] v3_1646635889_132;
   wire [1:0] itemTypeOut_w;
   wire [1:0] v3_1646635889_134;
   wire [1:0] v3_1646635889_135;
   wire [1:0] v3_1646635889_136;
   wire [1:0] v3_1646635889_137;
   wire [1:0] v3_1646635889_138;
   wire [1:0] v3_1646635889_139;
   wire [1:0] v3_1646635889_140;
   wire [1:0] v3_1646635889_141;
   wire [1:0] v3_1646635889_142;
   wire [1:0] v3_1646635889_143;
   wire [1:0] v3_1646635889_144;
   wire v3_1646635889_145;
   wire v3_1646635889_146;
   wire [1:0] v3_1646635889_147;
   wire [1:0] v3_1646635889_148;
   wire [1:0] v3_1646635889_149;
   wire [1:0] v3_1646635889_150;
   wire [1:0] v3_1646635889_151;
   wire [1:0] v3_1646635889_152;
   wire [1:0] v3_1646635889_153;
   wire [1:0] serviceTypeOut_w;
   wire [1:0] v3_1646635889_155;
   wire [1:0] v3_1646635889_156;
   wire [1:0] v3_1646635889_157;
   wire [1:0] v3_1646635889_158;
   wire [1:0] v3_1646635889_159;
   wire [1:0] v3_1646635889_160;
   wire [1:0] v3_1646635889_161;
   wire [1:0] v3_1646635889_162;
   wire [1:0] v3_1646635889_163;
   wire [1:0] v3_1646635889_164;
   wire [1:0] v3_1646635889_165;
   wire [1:0] v3_1646635889_166;
   wire [1:0] v3_1646635889_167;
   wire [1:0] v3_1646635889_168;
   wire [1:0] v3_1646635889_169;
   wire v3_1646635889_170;
   wire v3_1646635889_171;
   wire v3_1646635889_172;
   wire v3_1646635889_173;
   wire v3_1646635889_174;
   wire [7:0] v3_1646635889_175;
   wire [7:0] v3_1646635889_176;
   wire [7:0] inputValue_w;
   wire [7:0] v3_1646635889_178;
   wire [7:0] v3_1646635889_179;
   wire [7:0] v3_1646635889_180;
   wire [7:0] v3_1646635889_181;
   wire [7:0] v3_1646635889_182;
   wire [7:0] v3_1646635889_183;
   wire [7:0] v3_1646635889_184;
   wire [5:0] v3_1646635889_185;
   wire [7:0] v3_1646635889_186;
   wire [7:0] v3_1646635889_187;
   wire [7:0] v3_1646635889_188;
   wire [7:0] v3_1646635889_189;
   wire [7:0] v3_1646635889_190;
   wire [7:0] v3_1646635889_191;
   wire [7:0] v3_1646635889_192;
   wire [7:0] v3_1646635889_193;
   wire [7:0] v3_1646635889_194;
   wire [7:0] v3_1646635889_195;
   wire [7:0] v3_1646635889_196;
   wire [7:0] v3_1646635889_197;
   wire [7:0] v3_1646635889_198;
   wire [7:0] v3_1646635889_199;
   wire [7:0] v3_1646635889_200;
   wire [7:0] v3_1646635889_201;
   wire [7:0] v3_1646635889_202;
   wire [7:0] v3_1646635889_203;
   wire [7:0] v3_1646635889_204;
   wire [7:0] v3_1646635889_205;
   wire v3_1646635889_206;
   wire v3_1646635889_207;
   wire exchangeReady_w;
   wire v3_1646635889_209;
   wire v3_1646635889_210;
   wire v3_1646635889_211;
   wire v3_1646635889_212;
   wire v3_1646635889_213;
   wire v3_1646635889_214;
   wire v3_1646635889_215;
   wire v3_1646635889_216;
   wire v3_1646635889_217;
   wire v3_1646635889_218;
   wire v3_1646635889_219;
   wire [1:0] v3_1646635889_220;
   wire [1:0] v3_1646635889_221;
   wire [1:0] serviceCoinType_w;
   wire [1:0] v3_1646635889_223;
   wire [1:0] v3_1646635889_224;
   wire [1:0] v3_1646635889_225;
   wire [1:0] v3_1646635889_226;
   wire [1:0] v3_1646635889_227;
   wire [1:0] v3_1646635889_228;
   wire [1:0] v3_1646635889_229;
   wire [1:0] v3_1646635889_230;
   wire [1:0] v3_1646635889_231;
   wire [1:0] v3_1646635889_232;
   wire [1:0] v3_1646635889_233;
   wire [1:0] v3_1646635889_234;
   wire [1:0] v3_1646635889_235;
   wire [1:0] v3_1646635889_236;
   wire [1:0] v3_1646635889_237;
   wire [1:0] v3_1646635889_238;
   wire [1:0] v3_1646635889_239;
   wire [1:0] v3_1646635889_240;
   wire [1:0] v3_1646635889_241;
   wire [1:0] v3_1646635889_242;
   wire [1:0] v3_1646635889_243;
   wire [1:0] v3_1646635889_244;
   wire [1:0] v3_1646635889_245;
   wire [1:0] v3_1646635889_246;
   wire [1:0] v3_1646635889_247;
   wire [1:0] v3_1646635889_248;
   wire [7:0] v3_1646635889_249;
   wire [7:0] v3_1646635889_250;
   wire [7:0] serviceValue_w;
   wire [7:0] v3_1646635889_252;
   wire [7:0] v3_1646635889_253;
   wire [7:0] v3_1646635889_254;
   wire [7:0] v3_1646635889_255;
   wire [7:0] v3_1646635889_256;
   wire [7:0] v3_1646635889_257;
   wire [7:0] v3_1646635889_258;
   wire [7:0] v3_1646635889_259;
   wire [7:0] v3_1646635889_260;
   wire [7:0] v3_1646635889_261;
   wire [7:0] v3_1646635889_262;
   wire [7:0] v3_1646635889_263;
   wire [7:0] v3_1646635889_264;
   wire [7:0] v3_1646635889_265;
   wire [7:0] v3_1646635889_266;
   wire [7:0] v3_1646635889_267;
   wire [7:0] v3_1646635889_268;
   wire [7:0] v3_1646635889_269;
   wire [7:0] v3_1646635889_270;
   wire [7:0] v3_1646635889_271;
   wire [7:0] v3_1646635889_272;
   wire [7:0] v3_1646635889_273;
   wire [7:0] v3_1646635889_274;
   wire [7:0] v3_1646635889_275;
   wire [7:0] v3_1646635889_276;
   wire [7:0] v3_1646635889_277;
   wire [7:0] v3_1646635889_278;
   wire [7:0] v3_1646635889_279;
   wire [7:0] v3_1646635889_280;
   wire [7:0] v3_1646635889_281;
   wire [7:0] v3_1646635889_282;
   wire [7:0] v3_1646635889_283;
   wire v3_1646635889_284;
   wire [7:0] v3_1646635889_285;
   wire v3_1646635889_286;
   wire [7:0] v3_1646635889_287;
   wire v3_1646635889_288;
   wire [7:0] v3_1646635889_289;
   wire [7:0] v3_1646635889_290;
   wire [2:0] v3_1646635889_291;
   wire [2:0] v3_1646635889_292;
   wire [2:0] countNTD_50_w;
   wire [2:0] v3_1646635889_294;
   wire [2:0] v3_1646635889_295;
   wire [2:0] v3_1646635889_296;
   wire [2:0] v3_1646635889_297;
   wire [2:0] v3_1646635889_298;
   wire [2:0] v3_1646635889_299;
   wire [2:0] v3_1646635889_300;
   wire [2:0] v3_1646635889_301;
   wire [2:0] v3_1646635889_302;
   wire [2:0] v3_1646635889_303;
   wire [2:0] v3_1646635889_304;
   wire [2:0] v3_1646635889_305;
   wire [2:0] v3_1646635889_306;
   wire [2:0] v3_1646635889_307;
   wire [2:0] v3_1646635889_308;
   wire [2:0] v3_1646635889_309;
   wire [2:0] v3_1646635889_310;
   wire [2:0] v3_1646635889_311;
   wire [2:0] v3_1646635889_312;
   wire [2:0] v3_1646635889_313;
   wire [2:0] v3_1646635889_314;
   wire v3_1646635889_315;
   wire [3:0] v3_1646635889_316;
   wire [3:0] v3_1646635889_317;
   wire [3:0] v3_1646635889_318;
   wire [3:0] v3_1646635889_319;
   wire [3:0] v3_1646635889_320;
   wire [3:0] v3_1646635889_321;
   wire [3:0] v3_1646635889_322;
   wire [2:0] v3_1646635889_323;
   wire [2:0] v3_1646635889_324;
   wire [2:0] v3_1646635889_325;
   wire [2:0] v3_1646635889_326;
   wire [2:0] v3_1646635889_327;
   wire [2:0] countNTD_10_w;
   wire [2:0] v3_1646635889_329;
   wire [2:0] v3_1646635889_330;
   wire [2:0] v3_1646635889_331;
   wire [2:0] v3_1646635889_332;
   wire [2:0] v3_1646635889_333;
   wire [2:0] v3_1646635889_334;
   wire [2:0] v3_1646635889_335;
   wire [2:0] v3_1646635889_336;
   wire [2:0] v3_1646635889_337;
   wire [2:0] v3_1646635889_338;
   wire [2:0] v3_1646635889_339;
   wire [2:0] v3_1646635889_340;
   wire [2:0] v3_1646635889_341;
   wire [2:0] v3_1646635889_342;
   wire [2:0] v3_1646635889_343;
   wire [2:0] v3_1646635889_344;
   wire [2:0] v3_1646635889_345;
   wire [2:0] v3_1646635889_346;
   wire [2:0] v3_1646635889_347;
   wire [2:0] v3_1646635889_348;
   wire v3_1646635889_349;
   wire [3:0] v3_1646635889_350;
   wire [3:0] v3_1646635889_351;
   wire [3:0] v3_1646635889_352;
   wire [3:0] v3_1646635889_353;
   wire [3:0] v3_1646635889_354;
   wire [3:0] v3_1646635889_355;
   wire [2:0] v3_1646635889_356;
   wire [2:0] v3_1646635889_357;
   wire [2:0] v3_1646635889_358;
   wire [2:0] v3_1646635889_359;
   wire [2:0] countNTD_1_w;
   wire [2:0] v3_1646635889_361;
   wire [2:0] v3_1646635889_362;
   wire [2:0] v3_1646635889_363;
   wire [2:0] v3_1646635889_364;
   wire [2:0] v3_1646635889_365;
   wire [2:0] v3_1646635889_366;
   wire [2:0] v3_1646635889_367;
   wire [2:0] v3_1646635889_368;
   wire [2:0] v3_1646635889_369;
   wire [2:0] v3_1646635889_370;
   wire [2:0] v3_1646635889_371;
   wire [2:0] v3_1646635889_372;
   wire [2:0] v3_1646635889_373;
   wire [2:0] v3_1646635889_374;
   wire [2:0] v3_1646635889_375;
   wire [2:0] v3_1646635889_376;
   wire [2:0] v3_1646635889_377;
   wire [2:0] v3_1646635889_378;
   wire v3_1646635889_379;
   wire [3:0] v3_1646635889_380;
   wire [3:0] v3_1646635889_381;
   wire [3:0] v3_1646635889_382;
   wire [3:0] v3_1646635889_383;
   wire [3:0] v3_1646635889_384;
   wire [3:0] v3_1646635889_385;
   wire [2:0] v3_1646635889_386;
   wire [2:0] v3_1646635889_387;
   wire [2:0] v3_1646635889_388;
   wire [2:0] v3_1646635889_389;
   wire [2:0] countNTD_5_w;
   wire [2:0] v3_1646635889_391;
   wire [2:0] v3_1646635889_392;
   wire [2:0] v3_1646635889_393;
   wire [2:0] v3_1646635889_394;
   wire [2:0] v3_1646635889_395;
   wire [2:0] v3_1646635889_396;
   wire [2:0] v3_1646635889_397;
   wire [2:0] v3_1646635889_398;
   wire [2:0] v3_1646635889_399;
   wire [2:0] v3_1646635889_400;
   wire [2:0] v3_1646635889_401;
   wire [2:0] v3_1646635889_402;
   wire [2:0] v3_1646635889_403;
   wire [2:0] v3_1646635889_404;
   wire [2:0] v3_1646635889_405;
   wire [2:0] v3_1646635889_406;
   wire [2:0] v3_1646635889_407;
   wire [2:0] v3_1646635889_408;
   wire [2:0] v3_1646635889_409;
   wire [2:0] v3_1646635889_410;
   wire v3_1646635889_411;
   wire [3:0] v3_1646635889_412;
   wire [3:0] v3_1646635889_413;
   wire [3:0] v3_1646635889_414;
   wire [3:0] v3_1646635889_415;
   wire [3:0] v3_1646635889_416;
   wire [3:0] v3_1646635889_417;
   wire [2:0] v3_1646635889_418;
   wire [2:0] v3_1646635889_419;
   wire p;
   wire v3_1646635889_421;
   wire v3_1646635889_422;
   wire v3_1646635889_423;
   wire v3_1646635889_424;
   wire v3_1646635889_425;
   wire v3_1646635889_426;
   wire v3_1646635889_427;
   wire [7:0] outExchange;
   wire [7:0] v3_1646635889_429;
   wire [7:0] v3_1646635889_430;
   wire [7:0] v3_1646635889_431;
   wire [7:0] v3_1646635889_432;
   wire [4:0] v3_1646635889_433;
   wire [7:0] v3_1646635889_434;
   wire [7:0] v3_1646635889_435;
   wire [7:0] v3_1646635889_436;
   wire [7:0] v3_1646635889_437;
   wire [7:0] v3_1646635889_438;
   wire [7:0] v3_1646635889_439;
   wire [7:0] v3_1646635889_440;
   wire [7:0] v3_1646635889_441;
   wire [7:0] v3_1646635889_442;
   wire [7:0] v3_1646635889_443;
   wire [7:0] v3_1646635889_444;
   wire [7:0] v3_1646635889_445;
   wire [7:0] v3_1646635889_446;
   wire [7:0] v3_1646635889_447;
   wire [7:0] v3_1646635889_448;
   wire [7:0] v3_1646635889_449;
   wire [7:0] v3_1646635889_450;
   wire v3_1646635889_451;

   // Combinational Assignments
   assign id0 = 1'b0; 
   assign v3_1646635889_23 = v3_1646635889_62 ? v3_1646635889_61 : v3_1646635889_24;
   assign v3_1646635889_24 = coinOutNTD_50_w;
   assign coinOutNTD_50_w = v3_1646635889_60 ? v3_1646635889_56 : v3_1646635889_26;
   assign v3_1646635889_26 = v3_1646635889_55 ? v3_1646635889_54 : v3_1646635889_27;
   assign v3_1646635889_27 = v3_1646635889_53 ? v3_1646635889_32 : v3_1646635889_28;
   assign v3_1646635889_28 = v3_1646635889_51 ? v3_1646635889_43 : v3_1646635889_29;
   assign v3_1646635889_29 = v3_1646635889_41 ? v3_1646635889_32 : v3_1646635889_30;
   assign v3_1646635889_30 = v3_1646635889_39 ? v3_1646635889_32 : v3_1646635889_31;
   assign v3_1646635889_31 = v3_1646635889_37 ? v3_1646635889_33 : v3_1646635889_32;
   assign v3_1646635889_32 = coinOutNTD_50;
   assign v3_1646635889_33 = v3_1646635889_36 ? v3_1646635889_34 : v3_1646635889_32;
   assign v3_1646635889_34 = v3_1646635889_35;
   assign v3_1646635889_35 = 3'b000; 
   assign v3_1646635889_36 = countNTD_1 == v3_1646635889_35;
   assign v3_1646635889_37 = serviceValue >= v3_1646635889_38;
   assign v3_1646635889_38 = 8'b00000001; 
   assign v3_1646635889_39 = serviceCoinType == v3_1646635889_40;
   assign v3_1646635889_40 = 2'b10; 
   assign v3_1646635889_41 = serviceCoinType == v3_1646635889_42;
   assign v3_1646635889_42 = 2'b01; 
   assign v3_1646635889_43 = v3_1646635889_49 ? v3_1646635889_44 : v3_1646635889_32;
   assign v3_1646635889_44 = v3_1646635889_48 ? v3_1646635889_32 : v3_1646635889_45;
   assign v3_1646635889_45 = v3_1646635889_47;
   assign v3_1646635889_46 = 3'b001; 
   assign v3_1646635889_47 = coinOutNTD_50 + v3_1646635889_46;
   assign v3_1646635889_48 = countNTD_50 == v3_1646635889_35;
   assign v3_1646635889_49 = serviceValue >= v3_1646635889_50;
   assign v3_1646635889_50 = 8'b00110010; 
   assign v3_1646635889_51 = serviceCoinType == v3_1646635889_52;
   assign v3_1646635889_52 = 2'b00; 
   assign v3_1646635889_53 = ~exchangeReady;
   assign v3_1646635889_54 = v3_1646635889_35;
   assign v3_1646635889_55 = serviceTypeOut == v3_1646635889_52;
   assign v3_1646635889_56 = v3_1646635889_58 ? v3_1646635889_57 : v3_1646635889_32;
   assign v3_1646635889_57 = v3_1646635889_35;
   assign v3_1646635889_58 = ~v3_1646635889_59;
   assign v3_1646635889_59 = itemTypeIn == v3_1646635889_52;
   assign v3_1646635889_60 = serviceTypeOut == v3_1646635889_42;
   assign v3_1646635889_61 = v3_1646635889_35;
   assign v3_1646635889_62 = ~reset;
   assign v3_1646635889_63 = 3'b000; 
   assign v3_1646635889_64 = v3_1646635889_62 ? v3_1646635889_86 : v3_1646635889_65;
   assign v3_1646635889_65 = coinOutNTD_10_w;
   assign coinOutNTD_10_w = v3_1646635889_60 ? v3_1646635889_84 : v3_1646635889_67;
   assign v3_1646635889_67 = v3_1646635889_55 ? v3_1646635889_83 : v3_1646635889_68;
   assign v3_1646635889_68 = v3_1646635889_53 ? v3_1646635889_73 : v3_1646635889_69;
   assign v3_1646635889_69 = v3_1646635889_51 ? v3_1646635889_73 : v3_1646635889_70;
   assign v3_1646635889_70 = v3_1646635889_41 ? v3_1646635889_76 : v3_1646635889_71;
   assign v3_1646635889_71 = v3_1646635889_39 ? v3_1646635889_73 : v3_1646635889_72;
   assign v3_1646635889_72 = v3_1646635889_37 ? v3_1646635889_74 : v3_1646635889_73;
   assign v3_1646635889_73 = coinOutNTD_10;
   assign v3_1646635889_74 = v3_1646635889_36 ? v3_1646635889_75 : v3_1646635889_73;
   assign v3_1646635889_75 = v3_1646635889_35;
   assign v3_1646635889_76 = v3_1646635889_81 ? v3_1646635889_77 : v3_1646635889_73;
   assign v3_1646635889_77 = v3_1646635889_80 ? v3_1646635889_73 : v3_1646635889_78;
   assign v3_1646635889_78 = v3_1646635889_79;
   assign v3_1646635889_79 = coinOutNTD_10 + v3_1646635889_46;
   assign v3_1646635889_80 = countNTD_10 == v3_1646635889_35;
   assign v3_1646635889_81 = serviceValue >= v3_1646635889_82;
   assign v3_1646635889_82 = 8'b00001010; 
   assign v3_1646635889_83 = v3_1646635889_35;
   assign v3_1646635889_84 = v3_1646635889_58 ? v3_1646635889_85 : v3_1646635889_73;
   assign v3_1646635889_85 = v3_1646635889_35;
   assign v3_1646635889_86 = v3_1646635889_35;
   assign v3_1646635889_87 = 3'b000; 
   assign v3_1646635889_88 = v3_1646635889_62 ? v3_1646635889_110 : v3_1646635889_89;
   assign v3_1646635889_89 = coinOutNTD_5_w;
   assign coinOutNTD_5_w = v3_1646635889_60 ? v3_1646635889_108 : v3_1646635889_91;
   assign v3_1646635889_91 = v3_1646635889_55 ? v3_1646635889_107 : v3_1646635889_92;
   assign v3_1646635889_92 = v3_1646635889_53 ? v3_1646635889_97 : v3_1646635889_93;
   assign v3_1646635889_93 = v3_1646635889_51 ? v3_1646635889_97 : v3_1646635889_94;
   assign v3_1646635889_94 = v3_1646635889_41 ? v3_1646635889_97 : v3_1646635889_95;
   assign v3_1646635889_95 = v3_1646635889_39 ? v3_1646635889_100 : v3_1646635889_96;
   assign v3_1646635889_96 = v3_1646635889_37 ? v3_1646635889_98 : v3_1646635889_97;
   assign v3_1646635889_97 = coinOutNTD_5;
   assign v3_1646635889_98 = v3_1646635889_36 ? v3_1646635889_99 : v3_1646635889_97;
   assign v3_1646635889_99 = v3_1646635889_35;
   assign v3_1646635889_100 = v3_1646635889_105 ? v3_1646635889_101 : v3_1646635889_97;
   assign v3_1646635889_101 = v3_1646635889_104 ? v3_1646635889_97 : v3_1646635889_102;
   assign v3_1646635889_102 = v3_1646635889_103;
   assign v3_1646635889_103 = coinOutNTD_5 + v3_1646635889_46;
   assign v3_1646635889_104 = countNTD_5 == v3_1646635889_35;
   assign v3_1646635889_105 = serviceValue >= v3_1646635889_106;
   assign v3_1646635889_106 = 8'b00000101; 
   assign v3_1646635889_107 = v3_1646635889_35;
   assign v3_1646635889_108 = v3_1646635889_58 ? v3_1646635889_109 : v3_1646635889_97;
   assign v3_1646635889_109 = v3_1646635889_35;
   assign v3_1646635889_110 = v3_1646635889_35;
   assign v3_1646635889_111 = 3'b000; 
   assign v3_1646635889_112 = v3_1646635889_62 ? v3_1646635889_129 : v3_1646635889_113;
   assign v3_1646635889_113 = coinOutNTD_1_w;
   assign coinOutNTD_1_w = v3_1646635889_60 ? v3_1646635889_127 : v3_1646635889_115;
   assign v3_1646635889_115 = v3_1646635889_55 ? v3_1646635889_126 : v3_1646635889_116;
   assign v3_1646635889_116 = v3_1646635889_53 ? v3_1646635889_121 : v3_1646635889_117;
   assign v3_1646635889_117 = v3_1646635889_51 ? v3_1646635889_121 : v3_1646635889_118;
   assign v3_1646635889_118 = v3_1646635889_41 ? v3_1646635889_121 : v3_1646635889_119;
   assign v3_1646635889_119 = v3_1646635889_39 ? v3_1646635889_121 : v3_1646635889_120;
   assign v3_1646635889_120 = v3_1646635889_37 ? v3_1646635889_122 : v3_1646635889_121;
   assign v3_1646635889_121 = coinOutNTD_1;
   assign v3_1646635889_122 = v3_1646635889_36 ? v3_1646635889_125 : v3_1646635889_123;
   assign v3_1646635889_123 = v3_1646635889_124;
   assign v3_1646635889_124 = coinOutNTD_1 + v3_1646635889_46;
   assign v3_1646635889_125 = v3_1646635889_35;
   assign v3_1646635889_126 = v3_1646635889_35;
   assign v3_1646635889_127 = v3_1646635889_58 ? v3_1646635889_128 : v3_1646635889_121;
   assign v3_1646635889_128 = v3_1646635889_35;
   assign v3_1646635889_129 = v3_1646635889_35;
   assign v3_1646635889_130 = 3'b000; 
   assign v3_1646635889_131 = v3_1646635889_62 ? v3_1646635889_150 : v3_1646635889_132;
   assign v3_1646635889_132 = itemTypeOut_w;
   assign itemTypeOut_w = v3_1646635889_60 ? v3_1646635889_148 : v3_1646635889_134;
   assign v3_1646635889_134 = v3_1646635889_55 ? v3_1646635889_147 : v3_1646635889_135;
   assign v3_1646635889_135 = v3_1646635889_53 ? v3_1646635889_143 : v3_1646635889_136;
   assign v3_1646635889_136 = v3_1646635889_51 ? v3_1646635889_140 : v3_1646635889_137;
   assign v3_1646635889_137 = v3_1646635889_41 ? v3_1646635889_140 : v3_1646635889_138;
   assign v3_1646635889_138 = v3_1646635889_39 ? v3_1646635889_140 : v3_1646635889_139;
   assign v3_1646635889_139 = v3_1646635889_37 ? v3_1646635889_141 : v3_1646635889_140;
   assign v3_1646635889_140 = itemTypeOut;
   assign v3_1646635889_141 = v3_1646635889_36 ? v3_1646635889_142 : v3_1646635889_140;
   assign v3_1646635889_142 = v3_1646635889_52;
   assign v3_1646635889_143 = v3_1646635889_145 ? v3_1646635889_144 : v3_1646635889_140;
   assign v3_1646635889_144 = v3_1646635889_52;
   assign v3_1646635889_145 = ~v3_1646635889_146;
   assign v3_1646635889_146 = inputValue >= serviceValue;
   assign v3_1646635889_147 = v3_1646635889_52;
   assign v3_1646635889_148 = v3_1646635889_58 ? v3_1646635889_149 : v3_1646635889_140;
   assign v3_1646635889_149 = itemTypeIn;
   assign v3_1646635889_150 = v3_1646635889_52;
   assign v3_1646635889_151 = 2'b00; 
   assign v3_1646635889_152 = v3_1646635889_62 ? v3_1646635889_168 : v3_1646635889_153;
   assign v3_1646635889_153 = serviceTypeOut_w;
   assign serviceTypeOut_w = v3_1646635889_60 ? v3_1646635889_166 : v3_1646635889_155;
   assign v3_1646635889_155 = v3_1646635889_55 ? v3_1646635889_165 : v3_1646635889_156;
   assign v3_1646635889_156 = v3_1646635889_53 ? v3_1646635889_163 : v3_1646635889_157;
   assign v3_1646635889_157 = v3_1646635889_51 ? v3_1646635889_163 : v3_1646635889_158;
   assign v3_1646635889_158 = v3_1646635889_41 ? v3_1646635889_163 : v3_1646635889_159;
   assign v3_1646635889_159 = v3_1646635889_39 ? v3_1646635889_163 : v3_1646635889_160;
   assign v3_1646635889_160 = v3_1646635889_37 ? v3_1646635889_162 : v3_1646635889_161;
   assign v3_1646635889_161 = v3_1646635889_52;
   assign v3_1646635889_162 = v3_1646635889_36 ? v3_1646635889_164 : v3_1646635889_163;
   assign v3_1646635889_163 = serviceTypeOut;
   assign v3_1646635889_164 = v3_1646635889_52;
   assign v3_1646635889_165 = v3_1646635889_42;
   assign v3_1646635889_166 = v3_1646635889_58 ? v3_1646635889_167 : v3_1646635889_163;
   assign v3_1646635889_167 = v3_1646635889_40;
   assign v3_1646635889_168 = v3_1646635889_42;
   assign v3_1646635889_169 = 2'b00; 
   assign v3_1646635889_170 = v3_1646635889_62 ? v3_1646635889_172 : v3_1646635889_171;
   assign v3_1646635889_171 = initialized;
   assign v3_1646635889_172 = v3_1646635889_173;
   assign v3_1646635889_173 = 1'b1; 
   assign v3_1646635889_174 = 1'b0; 
   assign v3_1646635889_175 = v3_1646635889_62 ? v3_1646635889_203 : v3_1646635889_176;
   assign v3_1646635889_176 = inputValue_w;
   assign inputValue_w = v3_1646635889_60 ? v3_1646635889_179 : v3_1646635889_178;
   assign v3_1646635889_178 = inputValue;
   assign v3_1646635889_179 = v3_1646635889_58 ? v3_1646635889_180 : v3_1646635889_178;
   assign v3_1646635889_180 = v3_1646635889_202;
   assign v3_1646635889_181 = v3_1646635889_197;
   assign v3_1646635889_182 = v3_1646635889_192;
   assign v3_1646635889_183 = v3_1646635889_187;
   assign v3_1646635889_184 = v3_1646635889_186;
   assign v3_1646635889_185 = 6'b000000; 
   assign v3_1646635889_186 = {v3_1646635889_185, coinInNTD_50};
   assign v3_1646635889_187 = v3_1646635889_50 * v3_1646635889_184;
   assign v3_1646635889_188 = v3_1646635889_191;
   assign v3_1646635889_189 = v3_1646635889_190;
   assign v3_1646635889_190 = {v3_1646635889_185, coinInNTD_10};
   assign v3_1646635889_191 = v3_1646635889_82 * v3_1646635889_189;
   assign v3_1646635889_192 = v3_1646635889_183 + v3_1646635889_188;
   assign v3_1646635889_193 = v3_1646635889_196;
   assign v3_1646635889_194 = v3_1646635889_195;
   assign v3_1646635889_195 = {v3_1646635889_185, coinInNTD_5};
   assign v3_1646635889_196 = v3_1646635889_106 * v3_1646635889_194;
   assign v3_1646635889_197 = v3_1646635889_182 + v3_1646635889_193;
   assign v3_1646635889_198 = v3_1646635889_201;
   assign v3_1646635889_199 = v3_1646635889_200;
   assign v3_1646635889_200 = {v3_1646635889_185, coinInNTD_1};
   assign v3_1646635889_201 = v3_1646635889_38 * v3_1646635889_199;
   assign v3_1646635889_202 = v3_1646635889_181 + v3_1646635889_198;
   assign v3_1646635889_203 = v3_1646635889_204;
   assign v3_1646635889_204 = 8'b00000000; 
   assign v3_1646635889_205 = 8'b00000000; 
   assign v3_1646635889_206 = v3_1646635889_62 ? v3_1646635889_218 : v3_1646635889_207;
   assign v3_1646635889_207 = exchangeReady_w;
   assign exchangeReady_w = v3_1646635889_60 ? v3_1646635889_215 : v3_1646635889_209;
   assign v3_1646635889_209 = v3_1646635889_55 ? v3_1646635889_211 : v3_1646635889_210;
   assign v3_1646635889_210 = v3_1646635889_53 ? v3_1646635889_212 : v3_1646635889_211;
   assign v3_1646635889_211 = exchangeReady;
   assign v3_1646635889_212 = v3_1646635889_145 ? v3_1646635889_214 : v3_1646635889_213;
   assign v3_1646635889_213 = v3_1646635889_173;
   assign v3_1646635889_214 = v3_1646635889_173;
   assign v3_1646635889_215 = v3_1646635889_58 ? v3_1646635889_216 : v3_1646635889_211;
   assign v3_1646635889_216 = v3_1646635889_217;
   assign v3_1646635889_217 = 1'b0; 
   assign v3_1646635889_218 = v3_1646635889_217;
   assign v3_1646635889_219 = 1'b0; 
   assign v3_1646635889_220 = v3_1646635889_62 ? v3_1646635889_247 : v3_1646635889_221;
   assign v3_1646635889_221 = serviceCoinType_w;
   assign serviceCoinType_w = v3_1646635889_60 ? v3_1646635889_245 : v3_1646635889_223;
   assign v3_1646635889_223 = v3_1646635889_55 ? v3_1646635889_229 : v3_1646635889_224;
   assign v3_1646635889_224 = v3_1646635889_53 ? v3_1646635889_229 : v3_1646635889_225;
   assign v3_1646635889_225 = v3_1646635889_51 ? v3_1646635889_241 : v3_1646635889_226;
   assign v3_1646635889_226 = v3_1646635889_41 ? v3_1646635889_237 : v3_1646635889_227;
   assign v3_1646635889_227 = v3_1646635889_39 ? v3_1646635889_232 : v3_1646635889_228;
   assign v3_1646635889_228 = v3_1646635889_37 ? v3_1646635889_230 : v3_1646635889_229;
   assign v3_1646635889_229 = serviceCoinType;
   assign v3_1646635889_230 = v3_1646635889_36 ? v3_1646635889_231 : v3_1646635889_229;
   assign v3_1646635889_231 = v3_1646635889_52;
   assign v3_1646635889_232 = v3_1646635889_105 ? v3_1646635889_235 : v3_1646635889_233;
   assign v3_1646635889_233 = v3_1646635889_234;
   assign v3_1646635889_234 = 2'b11; 
   assign v3_1646635889_235 = v3_1646635889_104 ? v3_1646635889_236 : v3_1646635889_229;
   assign v3_1646635889_236 = v3_1646635889_234;
   assign v3_1646635889_237 = v3_1646635889_81 ? v3_1646635889_239 : v3_1646635889_238;
   assign v3_1646635889_238 = v3_1646635889_40;
   assign v3_1646635889_239 = v3_1646635889_80 ? v3_1646635889_240 : v3_1646635889_229;
   assign v3_1646635889_240 = v3_1646635889_40;
   assign v3_1646635889_241 = v3_1646635889_49 ? v3_1646635889_243 : v3_1646635889_242;
   assign v3_1646635889_242 = v3_1646635889_42;
   assign v3_1646635889_243 = v3_1646635889_48 ? v3_1646635889_244 : v3_1646635889_229;
   assign v3_1646635889_244 = v3_1646635889_42;
   assign v3_1646635889_245 = v3_1646635889_58 ? v3_1646635889_246 : v3_1646635889_229;
   assign v3_1646635889_246 = v3_1646635889_52;
   assign v3_1646635889_247 = v3_1646635889_52;
   assign v3_1646635889_248 = 2'b00; 
   assign v3_1646635889_249 = v3_1646635889_62 ? v3_1646635889_289 : v3_1646635889_250;
   assign v3_1646635889_250 = serviceValue_w;
   assign serviceValue_w = v3_1646635889_60 ? v3_1646635889_279 : v3_1646635889_252;
   assign v3_1646635889_252 = v3_1646635889_55 ? v3_1646635889_258 : v3_1646635889_253;
   assign v3_1646635889_253 = v3_1646635889_53 ? v3_1646635889_275 : v3_1646635889_254;
   assign v3_1646635889_254 = v3_1646635889_51 ? v3_1646635889_271 : v3_1646635889_255;
   assign v3_1646635889_255 = v3_1646635889_41 ? v3_1646635889_267 : v3_1646635889_256;
   assign v3_1646635889_256 = v3_1646635889_39 ? v3_1646635889_263 : v3_1646635889_257;
   assign v3_1646635889_257 = v3_1646635889_37 ? v3_1646635889_259 : v3_1646635889_258;
   assign v3_1646635889_258 = serviceValue;
   assign v3_1646635889_259 = v3_1646635889_36 ? v3_1646635889_262 : v3_1646635889_260;
   assign v3_1646635889_260 = v3_1646635889_261;
   assign v3_1646635889_261 = serviceValue - v3_1646635889_38;
   assign v3_1646635889_262 = inputValue;
   assign v3_1646635889_263 = v3_1646635889_105 ? v3_1646635889_264 : v3_1646635889_258;
   assign v3_1646635889_264 = v3_1646635889_104 ? v3_1646635889_258 : v3_1646635889_265;
   assign v3_1646635889_265 = v3_1646635889_266;
   assign v3_1646635889_266 = serviceValue - v3_1646635889_106;
   assign v3_1646635889_267 = v3_1646635889_81 ? v3_1646635889_268 : v3_1646635889_258;
   assign v3_1646635889_268 = v3_1646635889_80 ? v3_1646635889_258 : v3_1646635889_269;
   assign v3_1646635889_269 = v3_1646635889_270;
   assign v3_1646635889_270 = serviceValue - v3_1646635889_82;
   assign v3_1646635889_271 = v3_1646635889_49 ? v3_1646635889_272 : v3_1646635889_258;
   assign v3_1646635889_272 = v3_1646635889_48 ? v3_1646635889_258 : v3_1646635889_273;
   assign v3_1646635889_273 = v3_1646635889_274;
   assign v3_1646635889_274 = serviceValue - v3_1646635889_50;
   assign v3_1646635889_275 = v3_1646635889_145 ? v3_1646635889_278 : v3_1646635889_276;
   assign v3_1646635889_276 = v3_1646635889_277;
   assign v3_1646635889_277 = inputValue - serviceValue;
   assign v3_1646635889_278 = inputValue;
   assign v3_1646635889_279 = v3_1646635889_58 ? v3_1646635889_280 : v3_1646635889_258;
   assign v3_1646635889_280 = v3_1646635889_288 ? v3_1646635889_287 : v3_1646635889_281;
   assign v3_1646635889_281 = v3_1646635889_286 ? v3_1646635889_285 : v3_1646635889_282;
   assign v3_1646635889_282 = v3_1646635889_284 ? v3_1646635889_283 : v3_1646635889_204;
   assign v3_1646635889_283 = 8'b00010110; 
   assign v3_1646635889_284 = itemTypeIn == v3_1646635889_234;
   assign v3_1646635889_285 = 8'b00001111; 
   assign v3_1646635889_286 = itemTypeIn == v3_1646635889_40;
   assign v3_1646635889_287 = 8'b00001000; 
   assign v3_1646635889_288 = itemTypeIn == v3_1646635889_42;
   assign v3_1646635889_289 = v3_1646635889_204;
   assign v3_1646635889_290 = 8'b00000000; 
   assign v3_1646635889_291 = v3_1646635889_62 ? v3_1646635889_323 : v3_1646635889_292;
   assign v3_1646635889_292 = countNTD_50_w;
   assign countNTD_50_w = v3_1646635889_60 ? v3_1646635889_308 : v3_1646635889_294;
   assign v3_1646635889_294 = v3_1646635889_55 ? v3_1646635889_300 : v3_1646635889_295;
   assign v3_1646635889_295 = v3_1646635889_53 ? v3_1646635889_300 : v3_1646635889_296;
   assign v3_1646635889_296 = v3_1646635889_51 ? v3_1646635889_304 : v3_1646635889_297;
   assign v3_1646635889_297 = v3_1646635889_41 ? v3_1646635889_300 : v3_1646635889_298;
   assign v3_1646635889_298 = v3_1646635889_39 ? v3_1646635889_300 : v3_1646635889_299;
   assign v3_1646635889_299 = v3_1646635889_37 ? v3_1646635889_301 : v3_1646635889_300;
   assign v3_1646635889_300 = countNTD_50;
   assign v3_1646635889_301 = v3_1646635889_36 ? v3_1646635889_302 : v3_1646635889_300;
   assign v3_1646635889_302 = v3_1646635889_303;
   assign v3_1646635889_303 = countNTD_50 + coinOutNTD_50;
   assign v3_1646635889_304 = v3_1646635889_49 ? v3_1646635889_305 : v3_1646635889_300;
   assign v3_1646635889_305 = v3_1646635889_48 ? v3_1646635889_300 : v3_1646635889_306;
   assign v3_1646635889_306 = v3_1646635889_307;
   assign v3_1646635889_307 = countNTD_50 - v3_1646635889_46;
   assign v3_1646635889_308 = v3_1646635889_58 ? v3_1646635889_309 : v3_1646635889_300;
   assign v3_1646635889_309 = v3_1646635889_315 ? v3_1646635889_314 : v3_1646635889_310;
   assign v3_1646635889_310 = v3_1646635889_313;
   assign v3_1646635889_311 = v3_1646635889_312;
   assign v3_1646635889_312 = {v3_1646635889_217, coinInNTD_50};
   assign v3_1646635889_313 = countNTD_50 + v3_1646635889_311;
   assign v3_1646635889_314 = 3'b111; 
   assign v3_1646635889_315 = v3_1646635889_316 >= v3_1646635889_322;
   assign v3_1646635889_316 = v3_1646635889_321;
   assign v3_1646635889_317 = v3_1646635889_318;
   assign v3_1646635889_318 = {v3_1646635889_217, countNTD_50};
   assign v3_1646635889_319 = v3_1646635889_320;
   assign v3_1646635889_320 = {v3_1646635889_52, coinInNTD_50};
   assign v3_1646635889_321 = v3_1646635889_317 + v3_1646635889_319;
   assign v3_1646635889_322 = 4'b0111; 
   assign v3_1646635889_323 = v3_1646635889_324;
   assign v3_1646635889_324 = 3'b010; 
   assign v3_1646635889_325 = 3'b000; 
   assign v3_1646635889_326 = v3_1646635889_62 ? v3_1646635889_356 : v3_1646635889_327;
   assign v3_1646635889_327 = countNTD_10_w;
   assign countNTD_10_w = v3_1646635889_60 ? v3_1646635889_343 : v3_1646635889_329;
   assign v3_1646635889_329 = v3_1646635889_55 ? v3_1646635889_335 : v3_1646635889_330;
   assign v3_1646635889_330 = v3_1646635889_53 ? v3_1646635889_335 : v3_1646635889_331;
   assign v3_1646635889_331 = v3_1646635889_51 ? v3_1646635889_335 : v3_1646635889_332;
   assign v3_1646635889_332 = v3_1646635889_41 ? v3_1646635889_339 : v3_1646635889_333;
   assign v3_1646635889_333 = v3_1646635889_39 ? v3_1646635889_335 : v3_1646635889_334;
   assign v3_1646635889_334 = v3_1646635889_37 ? v3_1646635889_336 : v3_1646635889_335;
   assign v3_1646635889_335 = countNTD_10;
   assign v3_1646635889_336 = v3_1646635889_36 ? v3_1646635889_337 : v3_1646635889_335;
   assign v3_1646635889_337 = v3_1646635889_338;
   assign v3_1646635889_338 = countNTD_10 + coinOutNTD_10;
   assign v3_1646635889_339 = v3_1646635889_81 ? v3_1646635889_340 : v3_1646635889_335;
   assign v3_1646635889_340 = v3_1646635889_80 ? v3_1646635889_335 : v3_1646635889_341;
   assign v3_1646635889_341 = v3_1646635889_342;
   assign v3_1646635889_342 = countNTD_10 - v3_1646635889_46;
   assign v3_1646635889_343 = v3_1646635889_58 ? v3_1646635889_344 : v3_1646635889_335;
   assign v3_1646635889_344 = v3_1646635889_349 ? v3_1646635889_314 : v3_1646635889_345;
   assign v3_1646635889_345 = v3_1646635889_348;
   assign v3_1646635889_346 = v3_1646635889_347;
   assign v3_1646635889_347 = {v3_1646635889_217, coinInNTD_10};
   assign v3_1646635889_348 = countNTD_10 + v3_1646635889_346;
   assign v3_1646635889_349 = v3_1646635889_350 >= v3_1646635889_322;
   assign v3_1646635889_350 = v3_1646635889_355;
   assign v3_1646635889_351 = v3_1646635889_352;
   assign v3_1646635889_352 = {v3_1646635889_217, countNTD_10};
   assign v3_1646635889_353 = v3_1646635889_354;
   assign v3_1646635889_354 = {v3_1646635889_52, coinInNTD_10};
   assign v3_1646635889_355 = v3_1646635889_351 + v3_1646635889_353;
   assign v3_1646635889_356 = v3_1646635889_324;
   assign v3_1646635889_357 = 3'b000; 
   assign v3_1646635889_358 = v3_1646635889_62 ? v3_1646635889_386 : v3_1646635889_359;
   assign v3_1646635889_359 = countNTD_1_w;
   assign countNTD_1_w = v3_1646635889_60 ? v3_1646635889_373 : v3_1646635889_361;
   assign v3_1646635889_361 = v3_1646635889_55 ? v3_1646635889_367 : v3_1646635889_362;
   assign v3_1646635889_362 = v3_1646635889_53 ? v3_1646635889_367 : v3_1646635889_363;
   assign v3_1646635889_363 = v3_1646635889_51 ? v3_1646635889_367 : v3_1646635889_364;
   assign v3_1646635889_364 = v3_1646635889_41 ? v3_1646635889_367 : v3_1646635889_365;
   assign v3_1646635889_365 = v3_1646635889_39 ? v3_1646635889_367 : v3_1646635889_366;
   assign v3_1646635889_366 = v3_1646635889_37 ? v3_1646635889_368 : v3_1646635889_367;
   assign v3_1646635889_367 = countNTD_1;
   assign v3_1646635889_368 = v3_1646635889_36 ? v3_1646635889_371 : v3_1646635889_369;
   assign v3_1646635889_369 = v3_1646635889_370;
   assign v3_1646635889_370 = countNTD_1 - v3_1646635889_46;
   assign v3_1646635889_371 = v3_1646635889_372;
   assign v3_1646635889_372 = countNTD_1 + coinOutNTD_1;
   assign v3_1646635889_373 = v3_1646635889_58 ? v3_1646635889_374 : v3_1646635889_367;
   assign v3_1646635889_374 = v3_1646635889_379 ? v3_1646635889_314 : v3_1646635889_375;
   assign v3_1646635889_375 = v3_1646635889_378;
   assign v3_1646635889_376 = v3_1646635889_377;
   assign v3_1646635889_377 = {v3_1646635889_217, coinInNTD_1};
   assign v3_1646635889_378 = countNTD_1 + v3_1646635889_376;
   assign v3_1646635889_379 = v3_1646635889_380 >= v3_1646635889_322;
   assign v3_1646635889_380 = v3_1646635889_385;
   assign v3_1646635889_381 = v3_1646635889_382;
   assign v3_1646635889_382 = {v3_1646635889_217, countNTD_1};
   assign v3_1646635889_383 = v3_1646635889_384;
   assign v3_1646635889_384 = {v3_1646635889_52, coinInNTD_1};
   assign v3_1646635889_385 = v3_1646635889_381 + v3_1646635889_383;
   assign v3_1646635889_386 = v3_1646635889_324;
   assign v3_1646635889_387 = 3'b000; 
   assign v3_1646635889_388 = v3_1646635889_62 ? v3_1646635889_418 : v3_1646635889_389;
   assign v3_1646635889_389 = countNTD_5_w;
   assign countNTD_5_w = v3_1646635889_60 ? v3_1646635889_405 : v3_1646635889_391;
   assign v3_1646635889_391 = v3_1646635889_55 ? v3_1646635889_397 : v3_1646635889_392;
   assign v3_1646635889_392 = v3_1646635889_53 ? v3_1646635889_397 : v3_1646635889_393;
   assign v3_1646635889_393 = v3_1646635889_51 ? v3_1646635889_397 : v3_1646635889_394;
   assign v3_1646635889_394 = v3_1646635889_41 ? v3_1646635889_397 : v3_1646635889_395;
   assign v3_1646635889_395 = v3_1646635889_39 ? v3_1646635889_401 : v3_1646635889_396;
   assign v3_1646635889_396 = v3_1646635889_37 ? v3_1646635889_398 : v3_1646635889_397;
   assign v3_1646635889_397 = countNTD_5;
   assign v3_1646635889_398 = v3_1646635889_36 ? v3_1646635889_399 : v3_1646635889_397;
   assign v3_1646635889_399 = v3_1646635889_400;
   assign v3_1646635889_400 = countNTD_5 + coinOutNTD_5;
   assign v3_1646635889_401 = v3_1646635889_105 ? v3_1646635889_402 : v3_1646635889_397;
   assign v3_1646635889_402 = v3_1646635889_104 ? v3_1646635889_397 : v3_1646635889_403;
   assign v3_1646635889_403 = v3_1646635889_404;
   assign v3_1646635889_404 = countNTD_5 - v3_1646635889_46;
   assign v3_1646635889_405 = v3_1646635889_58 ? v3_1646635889_406 : v3_1646635889_397;
   assign v3_1646635889_406 = v3_1646635889_411 ? v3_1646635889_314 : v3_1646635889_407;
   assign v3_1646635889_407 = v3_1646635889_410;
   assign v3_1646635889_408 = v3_1646635889_409;
   assign v3_1646635889_409 = {v3_1646635889_217, coinInNTD_5};
   assign v3_1646635889_410 = countNTD_5 + v3_1646635889_408;
   assign v3_1646635889_411 = v3_1646635889_412 >= v3_1646635889_322;
   assign v3_1646635889_412 = v3_1646635889_417;
   assign v3_1646635889_413 = v3_1646635889_414;
   assign v3_1646635889_414 = {v3_1646635889_217, countNTD_5};
   assign v3_1646635889_415 = v3_1646635889_416;
   assign v3_1646635889_416 = {v3_1646635889_52, coinInNTD_5};
   assign v3_1646635889_417 = v3_1646635889_413 + v3_1646635889_415;
   assign v3_1646635889_418 = v3_1646635889_324;
   assign v3_1646635889_419 = 3'b000; 
   assign p = v3_1646635889_451;
   assign v3_1646635889_421 = v3_1646635889_425;
   assign v3_1646635889_422 = v3_1646635889_423;
   assign v3_1646635889_423 = initialized & v3_1646635889_55;
   assign v3_1646635889_424 = itemTypeOut == v3_1646635889_52;
   assign v3_1646635889_425 = v3_1646635889_422 & v3_1646635889_424;
   assign v3_1646635889_426 = ~v3_1646635889_427;
   assign v3_1646635889_427 = outExchange == inputValue;
   assign outExchange = v3_1646635889_450;
   assign v3_1646635889_429 = v3_1646635889_445;
   assign v3_1646635889_430 = v3_1646635889_440;
   assign v3_1646635889_431 = v3_1646635889_435;
   assign v3_1646635889_432 = v3_1646635889_434;
   assign v3_1646635889_433 = 5'b00000; 
   assign v3_1646635889_434 = {v3_1646635889_433, coinOutNTD_50};
   assign v3_1646635889_435 = v3_1646635889_50 * v3_1646635889_432;
   assign v3_1646635889_436 = v3_1646635889_439;
   assign v3_1646635889_437 = v3_1646635889_438;
   assign v3_1646635889_438 = {v3_1646635889_433, coinOutNTD_10};
   assign v3_1646635889_439 = v3_1646635889_82 * v3_1646635889_437;
   assign v3_1646635889_440 = v3_1646635889_431 + v3_1646635889_436;
   assign v3_1646635889_441 = v3_1646635889_444;
   assign v3_1646635889_442 = v3_1646635889_443;
   assign v3_1646635889_443 = {v3_1646635889_433, coinOutNTD_5};
   assign v3_1646635889_444 = v3_1646635889_106 * v3_1646635889_442;
   assign v3_1646635889_445 = v3_1646635889_430 + v3_1646635889_441;
   assign v3_1646635889_446 = v3_1646635889_449;
   assign v3_1646635889_447 = v3_1646635889_448;
   assign v3_1646635889_448 = {v3_1646635889_433, coinOutNTD_1};
   assign v3_1646635889_449 = v3_1646635889_38 * v3_1646635889_447;
   assign v3_1646635889_450 = v3_1646635889_429 + v3_1646635889_446;
   assign v3_1646635889_451 = v3_1646635889_421 & v3_1646635889_426;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      coinOutNTD_50 <= v3_1646635889_23;
      coinOutNTD_10 <= v3_1646635889_64;
      coinOutNTD_5 <= v3_1646635889_88;
      coinOutNTD_1 <= v3_1646635889_112;
      itemTypeOut <= v3_1646635889_131;
      serviceTypeOut <= v3_1646635889_152;
      initialized <= v3_1646635889_170;
      inputValue <= v3_1646635889_175;
      exchangeReady <= v3_1646635889_206;
      serviceCoinType <= v3_1646635889_220;
      serviceValue <= v3_1646635889_249;
      countNTD_50 <= v3_1646635889_291;
      countNTD_10 <= v3_1646635889_326;
      countNTD_1 <= v3_1646635889_358;
      countNTD_5 <= v3_1646635889_388;
   end
endmodule
